`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/19/2023 06:16:12 PM
// Design Name: 
// Module Name: sys_arr64
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module syst_arr64(
	input [15:0] inp_w0,inp_w64,inp_w128,inp_w192,inp_w256,inp_w320,inp_w384,inp_w448,inp_w512,inp_w576,inp_w640,inp_w704,inp_w768,inp_w832,inp_w896,inp_w960,inp_w1024,inp_w1088,inp_w1152,inp_w1216,inp_w1280,inp_w1344,inp_w1408,inp_w1472,inp_w1536,inp_w1600,inp_w1664,inp_w1728,inp_w1792,inp_w1856,inp_w1920,inp_w1984,inp_w2048,inp_w2112,inp_w2176,inp_w2240,inp_w2304,inp_w2368,inp_w2432,inp_w2496,inp_w2560,inp_w2624,inp_w2688,inp_w2752,inp_w2816,inp_w2880,inp_w2944,inp_w3008,inp_w3072,inp_w3136,inp_w3200,inp_w3264,inp_w3328,inp_w3392,inp_w3456,inp_w3520,inp_w3584,inp_w3648,inp_w3712,inp_w3776,inp_w3840,inp_w3904,inp_w3968,inp_w4032,inp_n0,inp_n1,inp_n2,inp_n3,inp_n4,inp_n5,inp_n6,inp_n7,inp_n8,inp_n9,inp_n10,inp_n11,inp_n12,inp_n13,inp_n14,inp_n15,inp_n16,inp_n17,inp_n18,inp_n19,inp_n20,inp_n21,inp_n22,inp_n23,inp_n24,inp_n25,inp_n26,inp_n27,inp_n28,inp_n29,inp_n30,inp_n31,inp_n32,inp_n33,inp_n34,inp_n35,inp_n36,inp_n37,inp_n38,inp_n39,inp_n40,inp_n41,inp_n42,inp_n43,inp_n44,inp_n45,inp_n46,inp_n47,inp_n48,inp_n49,inp_n50,inp_n51,inp_n52,inp_n53,inp_n54,inp_n55,inp_n56,inp_n57,inp_n58,inp_n59,inp_n60,inp_n61,inp_n62,inp_n63,
	output reg [15:0]  result_out0, result_out1, result_out2, result_out3, result_out4, result_out5, result_out6, result_out7, result_out8, result_out9, result_out10, result_out11, result_out12, result_out13, result_out14, result_out15, result_out16, result_out17, result_out18, result_out19, result_out20, result_out21, result_out22, result_out23, result_out24, result_out25, result_out26, result_out27, result_out28, result_out29, result_out30, result_out31, result_out32, result_out33, result_out34, result_out35, result_out36, result_out37, result_out38, result_out39, result_out40, result_out41, result_out42, result_out43, result_out44, result_out45, result_out46, result_out47, result_out48, result_out49, result_out50, result_out51, result_out52, result_out53, result_out54, result_out55, result_out56, result_out57, result_out58, result_out59, result_out60, result_out61, result_out62, result_out63,result_out64, result_out65, result_out66, result_out67, result_out68, result_out69, result_out70, result_out71, result_out72, result_out73, result_out74, result_out75, result_out76, result_out77, result_out78, result_out79, result_out80, result_out81, result_out82, result_out83, result_out84, result_out85, result_out86, result_out87, result_out88, result_out89, result_out90, result_out91, result_out92, result_out93, result_out94, result_out95, result_out96, result_out97, result_out98, result_out99, result_out100, result_out101, result_out102, result_out103, result_out104, result_out105, result_out106, result_out107, result_out108, result_out109, result_out110, result_out111, result_out112, result_out113, result_out114, result_out115, result_out116, result_out117, result_out118, result_out119, result_out120, result_out121, result_out122, result_out123, result_out124, result_out125, result_out126, result_out127, result_out128, result_out129, result_out130, result_out131, result_out132, result_out133, result_out134, result_out135, result_out136, result_out137, result_out138, result_out139, result_out140, result_out141, result_out142, result_out143, result_out144, result_out145, result_out146, result_out147, result_out148, result_out149, result_out150, result_out151, result_out152, result_out153, result_out154, result_out155, result_out156, result_out157, result_out158, result_out159, result_out160, result_out161, result_out162, result_out163, result_out164, result_out165, result_out166, result_out167, result_out168, result_out169, result_out170, result_out171, result_out172, result_out173, result_out174, result_out175, result_out176, result_out177, result_out178, result_out179, result_out180, result_out181, result_out182, result_out183, result_out184, result_out185, result_out186, result_out187, result_out188, result_out189, result_out190, result_out191, result_out192, result_out193, result_out194, result_out195, result_out196, result_out197, result_out198, result_out199, result_out200, result_out201, result_out202, result_out203, result_out204, result_out205, result_out206, result_out207, result_out208, result_out209, result_out210, result_out211, result_out212, result_out213, result_out214, result_out215, result_out216, result_out217, result_out218, result_out219, result_out220, result_out221, result_out222, result_out223, result_out224, result_out225, result_out226, result_out227, result_out228, result_out229, result_out230, result_out231, result_out232, result_out233, result_out234, result_out235, result_out236, result_out237, result_out238, result_out239, result_out240, result_out241, result_out242, result_out243, result_out244, result_out245, result_out246, result_out247, result_out248, result_out249, result_out250, result_out251, result_out252, result_out253, result_out254, result_out255, result_out256, result_out257, result_out258, result_out259, result_out260, result_out261, result_out262, result_out263, result_out264, result_out265, result_out266, result_out267, result_out268, result_out269, result_out270, result_out271, result_out272, result_out273, result_out274, result_out275, result_out276, result_out277, result_out278, result_out279, result_out280, result_out281, result_out282, result_out283, result_out284, result_out285, result_out286, result_out287, result_out288, result_out289, result_out290, result_out291, result_out292, result_out293, result_out294, result_out295, result_out296, result_out297, result_out298, result_out299, result_out300, result_out301, result_out302, result_out303, result_out304, result_out305, result_out306, result_out307, result_out308, result_out309, result_out310, result_out311, result_out312, result_out313, result_out314, result_out315, result_out316, result_out317, result_out318, result_out319, result_out320, result_out321, result_out322, result_out323, result_out324, result_out325, result_out326, result_out327, result_out328, result_out329, result_out330, result_out331, result_out332, result_out333, result_out334, result_out335, result_out336, result_out337, result_out338, result_out339, result_out340, result_out341, result_out342, result_out343, result_out344, result_out345, result_out346, result_out347, result_out348, result_out349, result_out350, result_out351, result_out352, result_out353, result_out354, result_out355, result_out356, result_out357, result_out358, result_out359, result_out360, result_out361, result_out362, result_out363, result_out364, result_out365, result_out366, result_out367, result_out368, result_out369, result_out370, result_out371, result_out372, result_out373, result_out374, result_out375, result_out376, result_out377, result_out378, result_out379, result_out380, result_out381, result_out382, result_out383, result_out384, result_out385, result_out386, result_out387, result_out388, result_out389, result_out390, result_out391, result_out392, result_out393, result_out394, result_out395, result_out396, result_out397, result_out398, result_out399, result_out400, result_out401, result_out402, result_out403, result_out404, result_out405, result_out406, result_out407, result_out408, result_out409, result_out410, result_out411, result_out412, result_out413, result_out414, result_out415, result_out416, result_out417, result_out418, result_out419, result_out420, result_out421, result_out422, result_out423, result_out424, result_out425, result_out426, result_out427, result_out428, result_out429, result_out430, result_out431, result_out432, result_out433, result_out434, result_out435, result_out436, result_out437, result_out438, result_out439, result_out440, result_out441, result_out442, result_out443, result_out444, result_out445, result_out446, result_out447, result_out448, result_out449, result_out450, result_out451, result_out452, result_out453, result_out454, result_out455, result_out456, result_out457, result_out458, result_out459, result_out460, result_out461, result_out462, result_out463, result_out464, result_out465, result_out466, result_out467, result_out468, result_out469, result_out470, result_out471, result_out472, result_out473, result_out474, result_out475, result_out476, result_out477, result_out478, result_out479, result_out480, result_out481, result_out482, result_out483, result_out484, result_out485, result_out486, result_out487, result_out488, result_out489, result_out490, result_out491, result_out492, result_out493, result_out494, result_out495, result_out496, result_out497, result_out498, result_out499, result_out500, result_out501, result_out502, result_out503, result_out504, result_out505, result_out506, result_out507, result_out508, result_out509, result_out510, result_out511, result_out512, result_out513, result_out514, result_out515, result_out516, result_out517, result_out518, result_out519, result_out520, result_out521, result_out522, result_out523, result_out524, result_out525, result_out526, result_out527, result_out528, result_out529, result_out530, result_out531, result_out532, result_out533, result_out534, result_out535, result_out536, result_out537, result_out538, result_out539, result_out540, result_out541, result_out542, result_out543, result_out544, result_out545, result_out546, result_out547, result_out548, result_out549, result_out550, result_out551, result_out552, result_out553, result_out554, result_out555, result_out556, result_out557, result_out558, result_out559, result_out560, result_out561, result_out562, result_out563, result_out564, result_out565, result_out566, result_out567, result_out568, result_out569, result_out570, result_out571, result_out572, result_out573, result_out574, result_out575, result_out576, result_out577, result_out578, result_out579, result_out580, result_out581, result_out582, result_out583, result_out584, result_out585, result_out586, result_out587, result_out588, result_out589, result_out590, result_out591, result_out592, result_out593, result_out594, result_out595, result_out596, result_out597, result_out598, result_out599, result_out600, result_out601, result_out602, result_out603, result_out604, result_out605, result_out606, result_out607, result_out608, result_out609, result_out610, result_out611, result_out612, result_out613, result_out614, result_out615, result_out616, result_out617, result_out618, result_out619, result_out620, result_out621, result_out622, result_out623, result_out624, result_out625, result_out626, result_out627, result_out628, result_out629, result_out630, result_out631, result_out632, result_out633, result_out634, result_out635, result_out636, result_out637, result_out638, result_out639, result_out640, result_out641, result_out642, result_out643, result_out644, result_out645, result_out646, result_out647, result_out648, result_out649, result_out650, result_out651, result_out652, result_out653, result_out654, result_out655, result_out656, result_out657, result_out658, result_out659, result_out660, result_out661, result_out662, result_out663, result_out664, result_out665, result_out666, result_out667, result_out668, result_out669, result_out670, result_out671, result_out672, result_out673, result_out674, result_out675, result_out676, result_out677, result_out678, result_out679, result_out680, result_out681, result_out682, result_out683, result_out684, result_out685, result_out686, result_out687, result_out688, result_out689, result_out690, result_out691, result_out692, result_out693, result_out694, result_out695, result_out696, result_out697, result_out698, result_out699, result_out700, result_out701, result_out702, result_out703, result_out704, result_out705, result_out706, result_out707, result_out708, result_out709, result_out710, result_out711, result_out712, result_out713, result_out714, result_out715, result_out716, result_out717, result_out718, result_out719, result_out720, result_out721, result_out722, result_out723, result_out724, result_out725, result_out726, result_out727, result_out728, result_out729, result_out730, result_out731, result_out732, result_out733, result_out734, result_out735, result_out736, result_out737, result_out738, result_out739, result_out740, result_out741, result_out742, result_out743, result_out744, result_out745, result_out746, result_out747, result_out748, result_out749, result_out750, result_out751, result_out752, result_out753, result_out754, result_out755, result_out756, result_out757, result_out758, result_out759, result_out760, result_out761, result_out762, result_out763, result_out764, result_out765, result_out766, result_out767, result_out768, result_out769, result_out770, result_out771, result_out772, result_out773, result_out774, result_out775, result_out776, result_out777, result_out778, result_out779, result_out780, result_out781, result_out782, result_out783, result_out784, result_out785, result_out786, result_out787, result_out788, result_out789, result_out790, result_out791, result_out792, result_out793, result_out794, result_out795, result_out796, result_out797, result_out798, result_out799, result_out800, result_out801, result_out802, result_out803, result_out804, result_out805, result_out806, result_out807, result_out808, result_out809, result_out810, result_out811, result_out812, result_out813, result_out814, result_out815, result_out816, result_out817, result_out818, result_out819, result_out820, result_out821, result_out822, result_out823, result_out824, result_out825, result_out826, result_out827, result_out828, result_out829, result_out830, result_out831, result_out832, result_out833, result_out834, result_out835, result_out836, result_out837, result_out838, result_out839, result_out840, result_out841, result_out842, result_out843, result_out844, result_out845, result_out846, result_out847, result_out848, result_out849, result_out850, result_out851, result_out852, result_out853, result_out854, result_out855, result_out856, result_out857, result_out858, result_out859, result_out860, result_out861, result_out862, result_out863, result_out864, result_out865, result_out866, result_out867, result_out868, result_out869, result_out870, result_out871, result_out872, result_out873, result_out874, result_out875, result_out876, result_out877, result_out878, result_out879, result_out880, result_out881, result_out882, result_out883, result_out884, result_out885, result_out886, result_out887, result_out888, result_out889, result_out890, result_out891, result_out892, result_out893, result_out894, result_out895, result_out896, result_out897, result_out898, result_out899, result_out900, result_out901, result_out902, result_out903, result_out904, result_out905, result_out906, result_out907, result_out908, result_out909, result_out910, result_out911, result_out912, result_out913, result_out914, result_out915, result_out916, result_out917, result_out918, result_out919, result_out920, result_out921, result_out922, result_out923, result_out924, result_out925, result_out926, result_out927, result_out928, result_out929, result_out930, result_out931, result_out932, result_out933, result_out934, result_out935, result_out936, result_out937, result_out938, result_out939, result_out940, result_out941, result_out942, result_out943, result_out944, result_out945, result_out946, result_out947, result_out948, result_out949, result_out950, result_out951, result_out952, result_out953, result_out954, result_out955, result_out956, result_out957, result_out958, result_out959, result_out960, result_out961, result_out962, result_out963, result_out964, result_out965, result_out966, result_out967, result_out968, result_out969, result_out970, result_out971, result_out972, result_out973, result_out974, result_out975, result_out976, result_out977, result_out978, result_out979, result_out980, result_out981, result_out982, result_out983, result_out984, result_out985, result_out986, result_out987, result_out988, result_out989, result_out990, result_out991, result_out992, result_out993, result_out994, result_out995, result_out996, result_out997, result_out998, result_out999, result_out1000, result_out1001, result_out1002, result_out1003, result_out1004, result_out1005, result_out1006, result_out1007, result_out1008, result_out1009, result_out1010, result_out1011, result_out1012, result_out1013, result_out1014, result_out1015, result_out1016, result_out1017, result_out1018, result_out1019, result_out1020, result_out1021, result_out1022, result_out1023, result_out1024, result_out1025, result_out1026, result_out1027, result_out1028, result_out1029, result_out1030, result_out1031, result_out1032, result_out1033, result_out1034, result_out1035, result_out1036, result_out1037, result_out1038, result_out1039, result_out1040, result_out1041, result_out1042, result_out1043, result_out1044, result_out1045, result_out1046, result_out1047, result_out1048, result_out1049, result_out1050, result_out1051, result_out1052, result_out1053, result_out1054, result_out1055, result_out1056, result_out1057, result_out1058, result_out1059, result_out1060, result_out1061, result_out1062, result_out1063, result_out1064, result_out1065, result_out1066, result_out1067, result_out1068, result_out1069, result_out1070, result_out1071, result_out1072, result_out1073, result_out1074, result_out1075, result_out1076, result_out1077, result_out1078, result_out1079, result_out1080, result_out1081, result_out1082, result_out1083, result_out1084, result_out1085, result_out1086, result_out1087, result_out1088, result_out1089, result_out1090, result_out1091, result_out1092, result_out1093, result_out1094, result_out1095, result_out1096, result_out1097, result_out1098, result_out1099, result_out1100, result_out1101, result_out1102, result_out1103, result_out1104, result_out1105, result_out1106, result_out1107, result_out1108, result_out1109, result_out1110, result_out1111, result_out1112, result_out1113, result_out1114, result_out1115, result_out1116, result_out1117, result_out1118, result_out1119, result_out1120, result_out1121, result_out1122, result_out1123, result_out1124, result_out1125, result_out1126, result_out1127, result_out1128, result_out1129, result_out1130, result_out1131, result_out1132, result_out1133, result_out1134, result_out1135, result_out1136, result_out1137, result_out1138, result_out1139, result_out1140, result_out1141, result_out1142, result_out1143, result_out1144, result_out1145, result_out1146, result_out1147, result_out1148, result_out1149, result_out1150, result_out1151, result_out1152, result_out1153, result_out1154, result_out1155, result_out1156, result_out1157, result_out1158, result_out1159, result_out1160, result_out1161, result_out1162, result_out1163, result_out1164, result_out1165, result_out1166, result_out1167, result_out1168, result_out1169, result_out1170, result_out1171, result_out1172, result_out1173, result_out1174, result_out1175, result_out1176, result_out1177, result_out1178, result_out1179, result_out1180, result_out1181, result_out1182, result_out1183, result_out1184, result_out1185, result_out1186, result_out1187, result_out1188, result_out1189, result_out1190, result_out1191, result_out1192, result_out1193, result_out1194, result_out1195, result_out1196, result_out1197, result_out1198, result_out1199, result_out1200, result_out1201, result_out1202, result_out1203, result_out1204, result_out1205, result_out1206, result_out1207, result_out1208, result_out1209, result_out1210, result_out1211, result_out1212, result_out1213, result_out1214, result_out1215, result_out1216, result_out1217, result_out1218, result_out1219, result_out1220, result_out1221, result_out1222, result_out1223, result_out1224, result_out1225, result_out1226, result_out1227, result_out1228, result_out1229, result_out1230, result_out1231, result_out1232, result_out1233, result_out1234, result_out1235, result_out1236, result_out1237, result_out1238, result_out1239, result_out1240, result_out1241, result_out1242, result_out1243, result_out1244, result_out1245, result_out1246, result_out1247, result_out1248, result_out1249, result_out1250, result_out1251, result_out1252, result_out1253, result_out1254, result_out1255, result_out1256, result_out1257, result_out1258, result_out1259, result_out1260, result_out1261, result_out1262, result_out1263, result_out1264, result_out1265, result_out1266, result_out1267, result_out1268, result_out1269, result_out1270, result_out1271, result_out1272, result_out1273, result_out1274, result_out1275, result_out1276, result_out1277, result_out1278, result_out1279, result_out1280, result_out1281, result_out1282, result_out1283, result_out1284, result_out1285, result_out1286, result_out1287, result_out1288, result_out1289, result_out1290, result_out1291, result_out1292, result_out1293, result_out1294, result_out1295, result_out1296, result_out1297, result_out1298, result_out1299, result_out1300, result_out1301, result_out1302, result_out1303, result_out1304, result_out1305, result_out1306, result_out1307, result_out1308, result_out1309, result_out1310, result_out1311, result_out1312, result_out1313, result_out1314, result_out1315, result_out1316, result_out1317, result_out1318, result_out1319, result_out1320, result_out1321, result_out1322, result_out1323, result_out1324, result_out1325, result_out1326, result_out1327, result_out1328, result_out1329, result_out1330, result_out1331, result_out1332, result_out1333, result_out1334, result_out1335, result_out1336, result_out1337, result_out1338, result_out1339, result_out1340, result_out1341, result_out1342, result_out1343, result_out1344, result_out1345, result_out1346, result_out1347, result_out1348, result_out1349, result_out1350, result_out1351, result_out1352, result_out1353, result_out1354, result_out1355, result_out1356, result_out1357, result_out1358, result_out1359, result_out1360, result_out1361, result_out1362, result_out1363, result_out1364, result_out1365, result_out1366, result_out1367, result_out1368, result_out1369, result_out1370, result_out1371, result_out1372, result_out1373, result_out1374, result_out1375, result_out1376, result_out1377, result_out1378, result_out1379, result_out1380, result_out1381, result_out1382, result_out1383, result_out1384, result_out1385, result_out1386, result_out1387, result_out1388, result_out1389, result_out1390, result_out1391, result_out1392, result_out1393, result_out1394, result_out1395, result_out1396, result_out1397, result_out1398, result_out1399, result_out1400, result_out1401, result_out1402, result_out1403, result_out1404, result_out1405, result_out1406, result_out1407, result_out1408, result_out1409, result_out1410, result_out1411, result_out1412, result_out1413, result_out1414, result_out1415, result_out1416, result_out1417, result_out1418, result_out1419, result_out1420, result_out1421, result_out1422, result_out1423, result_out1424, result_out1425, result_out1426, result_out1427, result_out1428, result_out1429, result_out1430, result_out1431, result_out1432, result_out1433, result_out1434, result_out1435, result_out1436, result_out1437, result_out1438, result_out1439, result_out1440, result_out1441, result_out1442, result_out1443, result_out1444, result_out1445, result_out1446, result_out1447, result_out1448, result_out1449, result_out1450, result_out1451, result_out1452, result_out1453, result_out1454, result_out1455, result_out1456, result_out1457, result_out1458, result_out1459, result_out1460, result_out1461, result_out1462, result_out1463, result_out1464, result_out1465, result_out1466, result_out1467, result_out1468, result_out1469, result_out1470, result_out1471, result_out1472, result_out1473, result_out1474, result_out1475, result_out1476, result_out1477, result_out1478, result_out1479, result_out1480, result_out1481, result_out1482, result_out1483, result_out1484, result_out1485, result_out1486, result_out1487, result_out1488, result_out1489, result_out1490, result_out1491, result_out1492, result_out1493, result_out1494, result_out1495, result_out1496, result_out1497, result_out1498, result_out1499, result_out1500, result_out1501, result_out1502, result_out1503, result_out1504, result_out1505, result_out1506, result_out1507, result_out1508, result_out1509, result_out1510, result_out1511, result_out1512, result_out1513, result_out1514, result_out1515, result_out1516, result_out1517, result_out1518, result_out1519, result_out1520, result_out1521, result_out1522, result_out1523, result_out1524, result_out1525, result_out1526, result_out1527, result_out1528, result_out1529, result_out1530, result_out1531, result_out1532, result_out1533, result_out1534, result_out1535, result_out1536, result_out1537, result_out1538, result_out1539, result_out1540, result_out1541, result_out1542, result_out1543, result_out1544, result_out1545, result_out1546, result_out1547, result_out1548, result_out1549, result_out1550, result_out1551, result_out1552, result_out1553, result_out1554, result_out1555, result_out1556, result_out1557, result_out1558, result_out1559, result_out1560, result_out1561, result_out1562, result_out1563, result_out1564, result_out1565, result_out1566, result_out1567, result_out1568, result_out1569, result_out1570, result_out1571, result_out1572, result_out1573, result_out1574, result_out1575, result_out1576, result_out1577, result_out1578, result_out1579, result_out1580, result_out1581, result_out1582, result_out1583, result_out1584, result_out1585, result_out1586, result_out1587, result_out1588, result_out1589, result_out1590, result_out1591, result_out1592, result_out1593, result_out1594, result_out1595, result_out1596, result_out1597, result_out1598, result_out1599, result_out1600, result_out1601, result_out1602, result_out1603, result_out1604, result_out1605, result_out1606, result_out1607, result_out1608, result_out1609, result_out1610, result_out1611, result_out1612, result_out1613, result_out1614, result_out1615, result_out1616, result_out1617, result_out1618, result_out1619, result_out1620, result_out1621, result_out1622, result_out1623, result_out1624, result_out1625, result_out1626, result_out1627, result_out1628, result_out1629, result_out1630, result_out1631, result_out1632, result_out1633, result_out1634, result_out1635, result_out1636, result_out1637, result_out1638, result_out1639, result_out1640, result_out1641, result_out1642, result_out1643, result_out1644, result_out1645, result_out1646, result_out1647, result_out1648, result_out1649, result_out1650, result_out1651, result_out1652, result_out1653, result_out1654, result_out1655, result_out1656, result_out1657, result_out1658, result_out1659, result_out1660, result_out1661, result_out1662, result_out1663, result_out1664, result_out1665, result_out1666, result_out1667, result_out1668, result_out1669, result_out1670, result_out1671, result_out1672, result_out1673, result_out1674, result_out1675, result_out1676, result_out1677, result_out1678, result_out1679, result_out1680, result_out1681, result_out1682, result_out1683, result_out1684, result_out1685, result_out1686, result_out1687, result_out1688, result_out1689, result_out1690, result_out1691, result_out1692, result_out1693, result_out1694, result_out1695, result_out1696, result_out1697, result_out1698, result_out1699, result_out1700, result_out1701, result_out1702, result_out1703, result_out1704, result_out1705, result_out1706, result_out1707, result_out1708, result_out1709, result_out1710, result_out1711, result_out1712, result_out1713, result_out1714, result_out1715, result_out1716, result_out1717, result_out1718, result_out1719, result_out1720, result_out1721, result_out1722, result_out1723, result_out1724, result_out1725, result_out1726, result_out1727, result_out1728, result_out1729, result_out1730, result_out1731, result_out1732, result_out1733, result_out1734, result_out1735, result_out1736, result_out1737, result_out1738, result_out1739, result_out1740, result_out1741, result_out1742, result_out1743, result_out1744, result_out1745, result_out1746, result_out1747, result_out1748, result_out1749, result_out1750, result_out1751, result_out1752, result_out1753, result_out1754, result_out1755, result_out1756, result_out1757, result_out1758, result_out1759, result_out1760, result_out1761, result_out1762, result_out1763, result_out1764, result_out1765, result_out1766, result_out1767, result_out1768, result_out1769, result_out1770, result_out1771, result_out1772, result_out1773, result_out1774, result_out1775, result_out1776, result_out1777, result_out1778, result_out1779, result_out1780, result_out1781, result_out1782, result_out1783, result_out1784, result_out1785, result_out1786, result_out1787, result_out1788, result_out1789, result_out1790, result_out1791, result_out1792, result_out1793, result_out1794, result_out1795, result_out1796, result_out1797, result_out1798, result_out1799, result_out1800, result_out1801, result_out1802, result_out1803, result_out1804, result_out1805, result_out1806, result_out1807, result_out1808, result_out1809, result_out1810, result_out1811, result_out1812, result_out1813, result_out1814, result_out1815, result_out1816, result_out1817, result_out1818, result_out1819, result_out1820, result_out1821, result_out1822, result_out1823, result_out1824, result_out1825, result_out1826, result_out1827, result_out1828, result_out1829, result_out1830, result_out1831, result_out1832, result_out1833, result_out1834, result_out1835, result_out1836, result_out1837, result_out1838, result_out1839, result_out1840, result_out1841, result_out1842, result_out1843, result_out1844, result_out1845, result_out1846, result_out1847, result_out1848, result_out1849, result_out1850, result_out1851, result_out1852, result_out1853, result_out1854, result_out1855, result_out1856, result_out1857, result_out1858, result_out1859, result_out1860, result_out1861, result_out1862, result_out1863, result_out1864, result_out1865, result_out1866, result_out1867, result_out1868, result_out1869, result_out1870, result_out1871, result_out1872, result_out1873, result_out1874, result_out1875, result_out1876, result_out1877, result_out1878, result_out1879, result_out1880, result_out1881, result_out1882, result_out1883, result_out1884, result_out1885, result_out1886, result_out1887, result_out1888, result_out1889, result_out1890, result_out1891, result_out1892, result_out1893, result_out1894, result_out1895, result_out1896, result_out1897, result_out1898, result_out1899, result_out1900, result_out1901, result_out1902, result_out1903, result_out1904, result_out1905, result_out1906, result_out1907, result_out1908, result_out1909, result_out1910, result_out1911, result_out1912, result_out1913, result_out1914, result_out1915, result_out1916, result_out1917, result_out1918, result_out1919, result_out1920, result_out1921, result_out1922, result_out1923, result_out1924, result_out1925, result_out1926, result_out1927, result_out1928, result_out1929, result_out1930, result_out1931, result_out1932, result_out1933, result_out1934, result_out1935, result_out1936, result_out1937, result_out1938, result_out1939, result_out1940, result_out1941, result_out1942, result_out1943, result_out1944, result_out1945, result_out1946, result_out1947, result_out1948, result_out1949, result_out1950, result_out1951, result_out1952, result_out1953, result_out1954, result_out1955, result_out1956, result_out1957, result_out1958, result_out1959, result_out1960, result_out1961, result_out1962, result_out1963, result_out1964, result_out1965, result_out1966, result_out1967, result_out1968, result_out1969, result_out1970, result_out1971, result_out1972, result_out1973, result_out1974, result_out1975, result_out1976, result_out1977, result_out1978, result_out1979, result_out1980, result_out1981, result_out1982, result_out1983, result_out1984, result_out1985, result_out1986, result_out1987, result_out1988, result_out1989, result_out1990, result_out1991, result_out1992, result_out1993, result_out1994, result_out1995, result_out1996, result_out1997, result_out1998, result_out1999, result_out2000, result_out2001, result_out2002, result_out2003, result_out2004, result_out2005, result_out2006, result_out2007, result_out2008, result_out2009, result_out2010, result_out2011, result_out2012, result_out2013, result_out2014, result_out2015, result_out2016, result_out2017, result_out2018, result_out2019, result_out2020, result_out2021, result_out2022, result_out2023, result_out2024, result_out2025, result_out2026, result_out2027, result_out2028, result_out2029, result_out2030, result_out2031, result_out2032, result_out2033, result_out2034, result_out2035, result_out2036, result_out2037, result_out2038, result_out2039, result_out2040, result_out2041, result_out2042, result_out2043, result_out2044, result_out2045, result_out2046, result_out2047, result_out2048, result_out2049, result_out2050, result_out2051, result_out2052, result_out2053, result_out2054, result_out2055, result_out2056, result_out2057, result_out2058, result_out2059, result_out2060, result_out2061, result_out2062, result_out2063, result_out2064, result_out2065, result_out2066, result_out2067, result_out2068, result_out2069, result_out2070, result_out2071, result_out2072, result_out2073, result_out2074, result_out2075, result_out2076, result_out2077, result_out2078, result_out2079, result_out2080, result_out2081, result_out2082, result_out2083, result_out2084, result_out2085, result_out2086, result_out2087, result_out2088, result_out2089, result_out2090, result_out2091, result_out2092, result_out2093, result_out2094, result_out2095, result_out2096, result_out2097, result_out2098, result_out2099, result_out2100, result_out2101, result_out2102, result_out2103, result_out2104, result_out2105, result_out2106, result_out2107, result_out2108, result_out2109, result_out2110, result_out2111, result_out2112, result_out2113, result_out2114, result_out2115, result_out2116, result_out2117, result_out2118, result_out2119, result_out2120, result_out2121, result_out2122, result_out2123, result_out2124, result_out2125, result_out2126, result_out2127, result_out2128, result_out2129, result_out2130, result_out2131, result_out2132, result_out2133, result_out2134, result_out2135, result_out2136, result_out2137, result_out2138, result_out2139, result_out2140, result_out2141, result_out2142, result_out2143, result_out2144, result_out2145, result_out2146, result_out2147, result_out2148, result_out2149, result_out2150, result_out2151, result_out2152, result_out2153, result_out2154, result_out2155, result_out2156, result_out2157, result_out2158, result_out2159, result_out2160, result_out2161, result_out2162, result_out2163, result_out2164, result_out2165, result_out2166, result_out2167, result_out2168, result_out2169, result_out2170, result_out2171, result_out2172, result_out2173, result_out2174, result_out2175, result_out2176, result_out2177, result_out2178, result_out2179, result_out2180, result_out2181, result_out2182, result_out2183, result_out2184, result_out2185, result_out2186, result_out2187, result_out2188, result_out2189, result_out2190, result_out2191, result_out2192, result_out2193, result_out2194, result_out2195, result_out2196, result_out2197, result_out2198, result_out2199, result_out2200, result_out2201, result_out2202, result_out2203, result_out2204, result_out2205, result_out2206, result_out2207, result_out2208, result_out2209, result_out2210, result_out2211, result_out2212, result_out2213, result_out2214, result_out2215, result_out2216, result_out2217, result_out2218, result_out2219, result_out2220, result_out2221, result_out2222, result_out2223, result_out2224, result_out2225, result_out2226, result_out2227, result_out2228, result_out2229, result_out2230, result_out2231, result_out2232, result_out2233, result_out2234, result_out2235, result_out2236, result_out2237, result_out2238, result_out2239, result_out2240, result_out2241, result_out2242, result_out2243, result_out2244, result_out2245, result_out2246, result_out2247, result_out2248, result_out2249, result_out2250, result_out2251, result_out2252, result_out2253, result_out2254, result_out2255, result_out2256, result_out2257, result_out2258, result_out2259, result_out2260, result_out2261, result_out2262, result_out2263, result_out2264, result_out2265, result_out2266, result_out2267, result_out2268, result_out2269, result_out2270, result_out2271, result_out2272, result_out2273, result_out2274, result_out2275, result_out2276, result_out2277, result_out2278, result_out2279, result_out2280, result_out2281, result_out2282, result_out2283, result_out2284, result_out2285, result_out2286, result_out2287, result_out2288, result_out2289, result_out2290, result_out2291, result_out2292, result_out2293, result_out2294, result_out2295, result_out2296, result_out2297, result_out2298, result_out2299, result_out2300, result_out2301, result_out2302, result_out2303, result_out2304, result_out2305, result_out2306, result_out2307, result_out2308, result_out2309, result_out2310, result_out2311, result_out2312, result_out2313, result_out2314, result_out2315, result_out2316, result_out2317, result_out2318, result_out2319, result_out2320, result_out2321, result_out2322, result_out2323, result_out2324, result_out2325, result_out2326, result_out2327, result_out2328, result_out2329, result_out2330, result_out2331, result_out2332, result_out2333, result_out2334, result_out2335, result_out2336, result_out2337, result_out2338, result_out2339, result_out2340, result_out2341, result_out2342, result_out2343, result_out2344, result_out2345, result_out2346, result_out2347, result_out2348, result_out2349, result_out2350, result_out2351, result_out2352, result_out2353, result_out2354, result_out2355, result_out2356, result_out2357, result_out2358, result_out2359, result_out2360, result_out2361, result_out2362, result_out2363, result_out2364, result_out2365, result_out2366, result_out2367, result_out2368, result_out2369, result_out2370, result_out2371, result_out2372, result_out2373, result_out2374, result_out2375, result_out2376, result_out2377, result_out2378, result_out2379, result_out2380, result_out2381, result_out2382, result_out2383, result_out2384, result_out2385, result_out2386, result_out2387, result_out2388, result_out2389, result_out2390, result_out2391, result_out2392, result_out2393, result_out2394, result_out2395, result_out2396, result_out2397, result_out2398, result_out2399, result_out2400, result_out2401, result_out2402, result_out2403, result_out2404, result_out2405, result_out2406, result_out2407, result_out2408, result_out2409, result_out2410, result_out2411, result_out2412, result_out2413, result_out2414, result_out2415, result_out2416, result_out2417, result_out2418, result_out2419, result_out2420, result_out2421, result_out2422, result_out2423, result_out2424, result_out2425, result_out2426, result_out2427, result_out2428, result_out2429, result_out2430, result_out2431, result_out2432, result_out2433, result_out2434, result_out2435, result_out2436, result_out2437, result_out2438, result_out2439, result_out2440, result_out2441, result_out2442, result_out2443, result_out2444, result_out2445, result_out2446, result_out2447, result_out2448, result_out2449, result_out2450, result_out2451, result_out2452, result_out2453, result_out2454, result_out2455, result_out2456, result_out2457, result_out2458, result_out2459, result_out2460, result_out2461, result_out2462, result_out2463, result_out2464, result_out2465, result_out2466, result_out2467, result_out2468, result_out2469, result_out2470, result_out2471, result_out2472, result_out2473, result_out2474, result_out2475, result_out2476, result_out2477, result_out2478, result_out2479, result_out2480, result_out2481, result_out2482, result_out2483, result_out2484, result_out2485, result_out2486, result_out2487, result_out2488, result_out2489, result_out2490, result_out2491, result_out2492, result_out2493, result_out2494, result_out2495, result_out2496, result_out2497, result_out2498, result_out2499, result_out2500, result_out2501, result_out2502, result_out2503, result_out2504, result_out2505, result_out2506, result_out2507, result_out2508, result_out2509, result_out2510, result_out2511, result_out2512, result_out2513, result_out2514, result_out2515, result_out2516, result_out2517, result_out2518, result_out2519, result_out2520, result_out2521, result_out2522, result_out2523, result_out2524, result_out2525, result_out2526, result_out2527, result_out2528, result_out2529, result_out2530, result_out2531, result_out2532, result_out2533, result_out2534, result_out2535, result_out2536, result_out2537, result_out2538, result_out2539, result_out2540, result_out2541, result_out2542, result_out2543, result_out2544, result_out2545, result_out2546, result_out2547, result_out2548, result_out2549, result_out2550, result_out2551, result_out2552, result_out2553, result_out2554, result_out2555, result_out2556, result_out2557, result_out2558, result_out2559, result_out2560, result_out2561, result_out2562, result_out2563, result_out2564, result_out2565, result_out2566, result_out2567, result_out2568, result_out2569, result_out2570, result_out2571, result_out2572, result_out2573, result_out2574, result_out2575, result_out2576, result_out2577, result_out2578, result_out2579, result_out2580, result_out2581, result_out2582, result_out2583, result_out2584, result_out2585, result_out2586, result_out2587, result_out2588, result_out2589, result_out2590, result_out2591, result_out2592, result_out2593, result_out2594, result_out2595, result_out2596, result_out2597, result_out2598, result_out2599, result_out2600, result_out2601, result_out2602, result_out2603, result_out2604, result_out2605, result_out2606, result_out2607, result_out2608, result_out2609, result_out2610, result_out2611, result_out2612, result_out2613, result_out2614, result_out2615, result_out2616, result_out2617, result_out2618, result_out2619, result_out2620, result_out2621, result_out2622, result_out2623, result_out2624, result_out2625, result_out2626, result_out2627, result_out2628, result_out2629, result_out2630, result_out2631, result_out2632, result_out2633, result_out2634, result_out2635, result_out2636, result_out2637, result_out2638, result_out2639, result_out2640, result_out2641, result_out2642, result_out2643, result_out2644, result_out2645, result_out2646, result_out2647, result_out2648, result_out2649, result_out2650, result_out2651, result_out2652, result_out2653, result_out2654, result_out2655, result_out2656, result_out2657, result_out2658, result_out2659, result_out2660, result_out2661, result_out2662, result_out2663, result_out2664, result_out2665, result_out2666, result_out2667, result_out2668, result_out2669, result_out2670, result_out2671, result_out2672, result_out2673, result_out2674, result_out2675, result_out2676, result_out2677, result_out2678, result_out2679, result_out2680, result_out2681, result_out2682, result_out2683, result_out2684, result_out2685, result_out2686, result_out2687, result_out2688, result_out2689, result_out2690, result_out2691, result_out2692, result_out2693, result_out2694, result_out2695, result_out2696, result_out2697, result_out2698, result_out2699, result_out2700, result_out2701, result_out2702, result_out2703, result_out2704, result_out2705, result_out2706, result_out2707, result_out2708, result_out2709, result_out2710, result_out2711, result_out2712, result_out2713, result_out2714, result_out2715, result_out2716, result_out2717, result_out2718, result_out2719, result_out2720, result_out2721, result_out2722, result_out2723, result_out2724, result_out2725, result_out2726, result_out2727, result_out2728, result_out2729, result_out2730, result_out2731, result_out2732, result_out2733, result_out2734, result_out2735, result_out2736, result_out2737, result_out2738, result_out2739, result_out2740, result_out2741, result_out2742, result_out2743, result_out2744, result_out2745, result_out2746, result_out2747, result_out2748, result_out2749, result_out2750, result_out2751, result_out2752, result_out2753, result_out2754, result_out2755, result_out2756, result_out2757, result_out2758, result_out2759, result_out2760, result_out2761, result_out2762, result_out2763, result_out2764, result_out2765, result_out2766, result_out2767, result_out2768, result_out2769, result_out2770, result_out2771, result_out2772, result_out2773, result_out2774, result_out2775, result_out2776, result_out2777, result_out2778, result_out2779, result_out2780, result_out2781, result_out2782, result_out2783, result_out2784, result_out2785, result_out2786, result_out2787, result_out2788, result_out2789, result_out2790, result_out2791, result_out2792, result_out2793, result_out2794, result_out2795, result_out2796, result_out2797, result_out2798, result_out2799, result_out2800, result_out2801, result_out2802, result_out2803, result_out2804, result_out2805, result_out2806, result_out2807, result_out2808, result_out2809, result_out2810, result_out2811, result_out2812, result_out2813, result_out2814, result_out2815, result_out2816, result_out2817, result_out2818, result_out2819, result_out2820, result_out2821, result_out2822, result_out2823, result_out2824, result_out2825, result_out2826, result_out2827, result_out2828, result_out2829, result_out2830, result_out2831, result_out2832, result_out2833, result_out2834, result_out2835, result_out2836, result_out2837, result_out2838, result_out2839, result_out2840, result_out2841, result_out2842, result_out2843, result_out2844, result_out2845, result_out2846, result_out2847, result_out2848, result_out2849, result_out2850, result_out2851, result_out2852, result_out2853, result_out2854, result_out2855, result_out2856, result_out2857, result_out2858, result_out2859, result_out2860, result_out2861, result_out2862, result_out2863, result_out2864, result_out2865, result_out2866, result_out2867, result_out2868, result_out2869, result_out2870, result_out2871, result_out2872, result_out2873, result_out2874, result_out2875, result_out2876, result_out2877, result_out2878, result_out2879, result_out2880, result_out2881, result_out2882, result_out2883, result_out2884, result_out2885, result_out2886, result_out2887, result_out2888, result_out2889, result_out2890, result_out2891, result_out2892, result_out2893, result_out2894, result_out2895, result_out2896, result_out2897, result_out2898, result_out2899, result_out2900, result_out2901, result_out2902, result_out2903, result_out2904, result_out2905, result_out2906, result_out2907, result_out2908, result_out2909, result_out2910, result_out2911, result_out2912, result_out2913, result_out2914, result_out2915, result_out2916, result_out2917, result_out2918, result_out2919, result_out2920, result_out2921, result_out2922, result_out2923, result_out2924, result_out2925, result_out2926, result_out2927, result_out2928, result_out2929, result_out2930, result_out2931, result_out2932, result_out2933, result_out2934, result_out2935, result_out2936, result_out2937, result_out2938, result_out2939, result_out2940, result_out2941, result_out2942, result_out2943, result_out2944, result_out2945, result_out2946, result_out2947, result_out2948, result_out2949, result_out2950, result_out2951, result_out2952, result_out2953, result_out2954, result_out2955, result_out2956, result_out2957, result_out2958, result_out2959, result_out2960, result_out2961, result_out2962, result_out2963, result_out2964, result_out2965, result_out2966, result_out2967, result_out2968, result_out2969, result_out2970, result_out2971, result_out2972, result_out2973, result_out2974, result_out2975, result_out2976, result_out2977, result_out2978, result_out2979, result_out2980, result_out2981, result_out2982, result_out2983, result_out2984, result_out2985, result_out2986, result_out2987, result_out2988, result_out2989, result_out2990, result_out2991, result_out2992, result_out2993, result_out2994, result_out2995, result_out2996, result_out2997, result_out2998, result_out2999, result_out3000, result_out3001, result_out3002, result_out3003, result_out3004, result_out3005, result_out3006, result_out3007, result_out3008, result_out3009, result_out3010, result_out3011, result_out3012, result_out3013, result_out3014, result_out3015, result_out3016, result_out3017, result_out3018, result_out3019, result_out3020, result_out3021, result_out3022, result_out3023, result_out3024, result_out3025, result_out3026, result_out3027, result_out3028, result_out3029, result_out3030, result_out3031, result_out3032, result_out3033, result_out3034, result_out3035, result_out3036, result_out3037, result_out3038, result_out3039, result_out3040, result_out3041, result_out3042, result_out3043, result_out3044, result_out3045, result_out3046, result_out3047, result_out3048, result_out3049, result_out3050, result_out3051, result_out3052, result_out3053, result_out3054, result_out3055, result_out3056, result_out3057, result_out3058, result_out3059, result_out3060, result_out3061, result_out3062, result_out3063, result_out3064, result_out3065, result_out3066, result_out3067, result_out3068, result_out3069, result_out3070, result_out3071, result_out3072, result_out3073, result_out3074, result_out3075, result_out3076, result_out3077, result_out3078, result_out3079, result_out3080, result_out3081, result_out3082, result_out3083, result_out3084, result_out3085, result_out3086, result_out3087, result_out3088, result_out3089, result_out3090, result_out3091, result_out3092, result_out3093, result_out3094, result_out3095, result_out3096, result_out3097, result_out3098, result_out3099, result_out3100, result_out3101, result_out3102, result_out3103, result_out3104, result_out3105, result_out3106, result_out3107, result_out3108, result_out3109, result_out3110, result_out3111, result_out3112, result_out3113, result_out3114, result_out3115, result_out3116, result_out3117, result_out3118, result_out3119, result_out3120, result_out3121, result_out3122, result_out3123, result_out3124, result_out3125, result_out3126, result_out3127, result_out3128, result_out3129, result_out3130, result_out3131, result_out3132, result_out3133, result_out3134, result_out3135, result_out3136, result_out3137, result_out3138, result_out3139, result_out3140, result_out3141, result_out3142, result_out3143, result_out3144, result_out3145, result_out3146, result_out3147, result_out3148, result_out3149, result_out3150, result_out3151, result_out3152, result_out3153, result_out3154, result_out3155, result_out3156, result_out3157, result_out3158, result_out3159, result_out3160, result_out3161, result_out3162, result_out3163, result_out3164, result_out3165, result_out3166, result_out3167, result_out3168, result_out3169, result_out3170, result_out3171, result_out3172, result_out3173, result_out3174, result_out3175, result_out3176, result_out3177, result_out3178, result_out3179, result_out3180, result_out3181, result_out3182, result_out3183, result_out3184, result_out3185, result_out3186, result_out3187, result_out3188, result_out3189, result_out3190, result_out3191, result_out3192, result_out3193, result_out3194, result_out3195, result_out3196, result_out3197, result_out3198, result_out3199, result_out3200, result_out3201, result_out3202, result_out3203, result_out3204, result_out3205, result_out3206, result_out3207, result_out3208, result_out3209, result_out3210, result_out3211, result_out3212, result_out3213, result_out3214, result_out3215, result_out3216, result_out3217, result_out3218, result_out3219, result_out3220, result_out3221, result_out3222, result_out3223, result_out3224, result_out3225, result_out3226, result_out3227, result_out3228, result_out3229, result_out3230, result_out3231, result_out3232, result_out3233, result_out3234, result_out3235, result_out3236, result_out3237, result_out3238, result_out3239, result_out3240, result_out3241, result_out3242, result_out3243, result_out3244, result_out3245, result_out3246, result_out3247, result_out3248, result_out3249, result_out3250, result_out3251, result_out3252, result_out3253, result_out3254, result_out3255, result_out3256, result_out3257, result_out3258, result_out3259, result_out3260, result_out3261, result_out3262, result_out3263, result_out3264, result_out3265, result_out3266, result_out3267, result_out3268, result_out3269, result_out3270, result_out3271, result_out3272, result_out3273, result_out3274, result_out3275, result_out3276, result_out3277, result_out3278, result_out3279, result_out3280, result_out3281, result_out3282, result_out3283, result_out3284, result_out3285, result_out3286, result_out3287, result_out3288, result_out3289, result_out3290, result_out3291, result_out3292, result_out3293, result_out3294, result_out3295, result_out3296, result_out3297, result_out3298, result_out3299, result_out3300, result_out3301, result_out3302, result_out3303, result_out3304, result_out3305, result_out3306, result_out3307, result_out3308, result_out3309, result_out3310, result_out3311, result_out3312, result_out3313, result_out3314, result_out3315, result_out3316, result_out3317, result_out3318, result_out3319, result_out3320, result_out3321, result_out3322, result_out3323, result_out3324, result_out3325, result_out3326, result_out3327, result_out3328, result_out3329, result_out3330, result_out3331, result_out3332, result_out3333, result_out3334, result_out3335, result_out3336, result_out3337, result_out3338, result_out3339, result_out3340, result_out3341, result_out3342, result_out3343, result_out3344, result_out3345, result_out3346, result_out3347, result_out3348, result_out3349, result_out3350, result_out3351, result_out3352, result_out3353, result_out3354, result_out3355, result_out3356, result_out3357, result_out3358, result_out3359, result_out3360, result_out3361, result_out3362, result_out3363, result_out3364, result_out3365, result_out3366, result_out3367, result_out3368, result_out3369, result_out3370, result_out3371, result_out3372, result_out3373, result_out3374, result_out3375, result_out3376, result_out3377, result_out3378, result_out3379, result_out3380, result_out3381, result_out3382, result_out3383, result_out3384, result_out3385, result_out3386, result_out3387, result_out3388, result_out3389, result_out3390, result_out3391, result_out3392, result_out3393, result_out3394, result_out3395, result_out3396, result_out3397, result_out3398, result_out3399, result_out3400, result_out3401, result_out3402, result_out3403, result_out3404, result_out3405, result_out3406, result_out3407, result_out3408, result_out3409, result_out3410, result_out3411, result_out3412, result_out3413, result_out3414, result_out3415, result_out3416, result_out3417, result_out3418, result_out3419, result_out3420, result_out3421, result_out3422, result_out3423, result_out3424, result_out3425, result_out3426, result_out3427, result_out3428, result_out3429, result_out3430, result_out3431, result_out3432, result_out3433, result_out3434, result_out3435, result_out3436, result_out3437, result_out3438, result_out3439, result_out3440, result_out3441, result_out3442, result_out3443, result_out3444, result_out3445, result_out3446, result_out3447, result_out3448, result_out3449, result_out3450, result_out3451, result_out3452, result_out3453, result_out3454, result_out3455, result_out3456, result_out3457, result_out3458, result_out3459, result_out3460, result_out3461, result_out3462, result_out3463, result_out3464, result_out3465, result_out3466, result_out3467, result_out3468, result_out3469, result_out3470, result_out3471, result_out3472, result_out3473, result_out3474, result_out3475, result_out3476, result_out3477, result_out3478, result_out3479, result_out3480, result_out3481, result_out3482, result_out3483, result_out3484, result_out3485, result_out3486, result_out3487, result_out3488, result_out3489, result_out3490, result_out3491, result_out3492, result_out3493, result_out3494, result_out3495, result_out3496, result_out3497, result_out3498, result_out3499, result_out3500, result_out3501, result_out3502, result_out3503, result_out3504, result_out3505, result_out3506, result_out3507, result_out3508, result_out3509, result_out3510, result_out3511, result_out3512, result_out3513, result_out3514, result_out3515, result_out3516, result_out3517, result_out3518, result_out3519, result_out3520, result_out3521, result_out3522, result_out3523, result_out3524, result_out3525, result_out3526, result_out3527, result_out3528, result_out3529, result_out3530, result_out3531, result_out3532, result_out3533, result_out3534, result_out3535, result_out3536, result_out3537, result_out3538, result_out3539, result_out3540, result_out3541, result_out3542, result_out3543, result_out3544, result_out3545, result_out3546, result_out3547, result_out3548, result_out3549, result_out3550, result_out3551, result_out3552, result_out3553, result_out3554, result_out3555, result_out3556, result_out3557, result_out3558, result_out3559, result_out3560, result_out3561, result_out3562, result_out3563, result_out3564, result_out3565, result_out3566, result_out3567, result_out3568, result_out3569, result_out3570, result_out3571, result_out3572, result_out3573, result_out3574, result_out3575, result_out3576, result_out3577, result_out3578, result_out3579, result_out3580, result_out3581, result_out3582, result_out3583, result_out3584, result_out3585, result_out3586, result_out3587, result_out3588, result_out3589, result_out3590, result_out3591, result_out3592, result_out3593, result_out3594, result_out3595, result_out3596, result_out3597, result_out3598, result_out3599, result_out3600, result_out3601, result_out3602, result_out3603, result_out3604, result_out3605, result_out3606, result_out3607, result_out3608, result_out3609, result_out3610, result_out3611, result_out3612, result_out3613, result_out3614, result_out3615, result_out3616, result_out3617, result_out3618, result_out3619, result_out3620, result_out3621, result_out3622, result_out3623, result_out3624, result_out3625, result_out3626, result_out3627, result_out3628, result_out3629, result_out3630, result_out3631, result_out3632, result_out3633, result_out3634, result_out3635, result_out3636, result_out3637, result_out3638, result_out3639, result_out3640, result_out3641, result_out3642, result_out3643, result_out3644, result_out3645, result_out3646, result_out3647, result_out3648, result_out3649, result_out3650, result_out3651, result_out3652, result_out3653, result_out3654, result_out3655, result_out3656, result_out3657, result_out3658, result_out3659, result_out3660, result_out3661, result_out3662, result_out3663, result_out3664, result_out3665, result_out3666, result_out3667, result_out3668, result_out3669, result_out3670, result_out3671, result_out3672, result_out3673, result_out3674, result_out3675, result_out3676, result_out3677, result_out3678, result_out3679, result_out3680, result_out3681, result_out3682, result_out3683, result_out3684, result_out3685, result_out3686, result_out3687, result_out3688, result_out3689, result_out3690, result_out3691, result_out3692, result_out3693, result_out3694, result_out3695, result_out3696, result_out3697, result_out3698, result_out3699, result_out3700, result_out3701, result_out3702, result_out3703, result_out3704, result_out3705, result_out3706, result_out3707, result_out3708, result_out3709, result_out3710, result_out3711, result_out3712, result_out3713, result_out3714, result_out3715, result_out3716, result_out3717, result_out3718, result_out3719, result_out3720, result_out3721, result_out3722, result_out3723, result_out3724, result_out3725, result_out3726, result_out3727, result_out3728, result_out3729, result_out3730, result_out3731, result_out3732, result_out3733, result_out3734, result_out3735, result_out3736, result_out3737, result_out3738, result_out3739, result_out3740, result_out3741, result_out3742, result_out3743, result_out3744, result_out3745, result_out3746, result_out3747, result_out3748, result_out3749, result_out3750, result_out3751, result_out3752, result_out3753, result_out3754, result_out3755, result_out3756, result_out3757, result_out3758, result_out3759, result_out3760, result_out3761, result_out3762, result_out3763, result_out3764, result_out3765, result_out3766, result_out3767, result_out3768, result_out3769, result_out3770, result_out3771, result_out3772, result_out3773, result_out3774, result_out3775, result_out3776, result_out3777, result_out3778, result_out3779, result_out3780, result_out3781, result_out3782, result_out3783, result_out3784, result_out3785, result_out3786, result_out3787, result_out3788, result_out3789, result_out3790, result_out3791, result_out3792, result_out3793, result_out3794, result_out3795, result_out3796, result_out3797, result_out3798, result_out3799, result_out3800, result_out3801, result_out3802, result_out3803, result_out3804, result_out3805, result_out3806, result_out3807, result_out3808, result_out3809, result_out3810, result_out3811, result_out3812, result_out3813, result_out3814, result_out3815, result_out3816, result_out3817, result_out3818, result_out3819, result_out3820, result_out3821, result_out3822, result_out3823, result_out3824, result_out3825, result_out3826, result_out3827, result_out3828, result_out3829, result_out3830, result_out3831, result_out3832, result_out3833, result_out3834, result_out3835, result_out3836, result_out3837, result_out3838, result_out3839, result_out3840, result_out3841, result_out3842, result_out3843, result_out3844, result_out3845, result_out3846, result_out3847, result_out3848, result_out3849, result_out3850, result_out3851, result_out3852, result_out3853, result_out3854, result_out3855, result_out3856, result_out3857, result_out3858, result_out3859, result_out3860, result_out3861, result_out3862, result_out3863, result_out3864, result_out3865, result_out3866, result_out3867, result_out3868, result_out3869, result_out3870, result_out3871, result_out3872, result_out3873, result_out3874, result_out3875, result_out3876, result_out3877, result_out3878, result_out3879, result_out3880, result_out3881, result_out3882, result_out3883, result_out3884, result_out3885, result_out3886, result_out3887, result_out3888, result_out3889, result_out3890, result_out3891, result_out3892, result_out3893, result_out3894, result_out3895, result_out3896, result_out3897, result_out3898, result_out3899, result_out3900, result_out3901, result_out3902, result_out3903, result_out3904, result_out3905, result_out3906, result_out3907, result_out3908, result_out3909, result_out3910, result_out3911, result_out3912, result_out3913, result_out3914, result_out3915, result_out3916, result_out3917, result_out3918, result_out3919, result_out3920, result_out3921, result_out3922, result_out3923, result_out3924, result_out3925, result_out3926, result_out3927, result_out3928, result_out3929, result_out3930, result_out3931, result_out3932, result_out3933, result_out3934, result_out3935, result_out3936, result_out3937, result_out3938, result_out3939, result_out3940, result_out3941, result_out3942, result_out3943, result_out3944, result_out3945, result_out3946, result_out3947, result_out3948, result_out3949, result_out3950, result_out3951, result_out3952, result_out3953, result_out3954, result_out3955, result_out3956, result_out3957, result_out3958, result_out3959, result_out3960, result_out3961, result_out3962, result_out3963, result_out3964, result_out3965, result_out3966, result_out3967, result_out3968, result_out3969, result_out3970, result_out3971, result_out3972, result_out3973, result_out3974, result_out3975, result_out3976, result_out3977, result_out3978, result_out3979, result_out3980, result_out3981, result_out3982, result_out3983, result_out3984, result_out3985, result_out3986, result_out3987, result_out3988, result_out3989, result_out3990, result_out3991, result_out3992, result_out3993, result_out3994, result_out3995, result_out3996, result_out3997, result_out3998, result_out3999, result_out4000, result_out4001, result_out4002, result_out4003, result_out4004, result_out4005, result_out4006, result_out4007, result_out4008, result_out4009, result_out4010, result_out4011, result_out4012, result_out4013, result_out4014, result_out4015, result_out4016, result_out4017, result_out4018, result_out4019, result_out4020, result_out4021, result_out4022, result_out4023, result_out4024, result_out4025, result_out4026, result_out4027, result_out4028, result_out4029, result_out4030, result_out4031, result_out4032, result_out4033, result_out4034, result_out4035, result_out4036, result_out4037, result_out4038, result_out4039, result_out4040, result_out4041, result_out4042, result_out4043, result_out4044, result_out4045, result_out4046, result_out4047, result_out4048, result_out4049, result_out4050, result_out4051, result_out4052, result_out4053, result_out4054, result_out4055, result_out4056, result_out4057, result_out4058, result_out4059, result_out4060, result_out4061, result_out4062, result_out4063, result_out4064, result_out4065, result_out4066, result_out4067, result_out4068, result_out4069, result_out4070, result_out4071, result_out4072, result_out4073, result_out4074, result_out4075, result_out4076, result_out4077, result_out4078, result_out4079, result_out4080, result_out4081, result_out4082, result_out4083, result_out4084, result_out4085, result_out4086, result_out4087, result_out4088, result_out4089, result_out4090, result_out4091, result_out4092, result_out4093, result_out4094, result_out4095, 
	output reg done,
	input clk,rst
); 

reg [7:0] count;

wire  [15:0] out_s0;
wire  [15:0] out_s1;
wire  [15:0] out_s2;
wire  [15:0] out_s3;
wire  [15:0] out_s4;
wire  [15:0] out_s5;
wire  [15:0] out_s6;
wire  [15:0] out_s7;
wire  [15:0] out_s8;
wire  [15:0] out_s9;
wire  [15:0] out_s10;
wire  [15:0] out_s11;
wire  [15:0] out_s12;
wire  [15:0] out_s13;
wire  [15:0] out_s14;
wire  [15:0] out_s15;
wire  [15:0] out_s16;
wire  [15:0] out_s17;
wire  [15:0] out_s18;
wire  [15:0] out_s19;
wire  [15:0] out_s20;
wire  [15:0] out_s21;
wire  [15:0] out_s22;
wire  [15:0] out_s23;
wire  [15:0] out_s24;
wire  [15:0] out_s25;
wire  [15:0] out_s26;
wire  [15:0] out_s27;
wire  [15:0] out_s28;
wire  [15:0] out_s29;
wire  [15:0] out_s30;
wire  [15:0] out_s31;
wire  [15:0] out_s32;
wire  [15:0] out_s33;
wire  [15:0] out_s34;
wire  [15:0] out_s35;
wire  [15:0] out_s36;
wire  [15:0] out_s37;
wire  [15:0] out_s38;
wire  [15:0] out_s39;
wire  [15:0] out_s40;
wire  [15:0] out_s41;
wire  [15:0] out_s42;
wire  [15:0] out_s43;
wire  [15:0] out_s44;
wire  [15:0] out_s45;
wire  [15:0] out_s46;
wire  [15:0] out_s47;
wire  [15:0] out_s48;
wire  [15:0] out_s49;
wire  [15:0] out_s50;
wire  [15:0] out_s51;
wire  [15:0] out_s52;
wire  [15:0] out_s53;
wire  [15:0] out_s54;
wire  [15:0] out_s55;
wire  [15:0] out_s56;
wire  [15:0] out_s57;
wire  [15:0] out_s58;
wire  [15:0] out_s59;
wire  [15:0] out_s60;
wire  [15:0] out_s61;
wire  [15:0] out_s62;
wire  [15:0] out_s63;
wire  [15:0] out_s64;
wire  [15:0] out_s65;
wire  [15:0] out_s66;
wire  [15:0] out_s67;
wire  [15:0] out_s68;
wire  [15:0] out_s69;
wire  [15:0] out_s70;
wire  [15:0] out_s71;
wire  [15:0] out_s72;
wire  [15:0] out_s73;
wire  [15:0] out_s74;
wire  [15:0] out_s75;
wire  [15:0] out_s76;
wire  [15:0] out_s77;
wire  [15:0] out_s78;
wire  [15:0] out_s79;
wire  [15:0] out_s80;
wire  [15:0] out_s81;
wire  [15:0] out_s82;
wire  [15:0] out_s83;
wire  [15:0] out_s84;
wire  [15:0] out_s85;
wire  [15:0] out_s86;
wire  [15:0] out_s87;
wire  [15:0] out_s88;
wire  [15:0] out_s89;
wire  [15:0] out_s90;
wire  [15:0] out_s91;
wire  [15:0] out_s92;
wire  [15:0] out_s93;
wire  [15:0] out_s94;
wire  [15:0] out_s95;
wire  [15:0] out_s96;
wire  [15:0] out_s97;
wire  [15:0] out_s98;
wire  [15:0] out_s99;
wire  [15:0] out_s100;
wire  [15:0] out_s101;
wire  [15:0] out_s102;
wire  [15:0] out_s103;
wire  [15:0] out_s104;
wire  [15:0] out_s105;
wire  [15:0] out_s106;
wire  [15:0] out_s107;
wire  [15:0] out_s108;
wire  [15:0] out_s109;
wire  [15:0] out_s110;
wire  [15:0] out_s111;
wire  [15:0] out_s112;
wire  [15:0] out_s113;
wire  [15:0] out_s114;
wire  [15:0] out_s115;
wire  [15:0] out_s116;
wire  [15:0] out_s117;
wire  [15:0] out_s118;
wire  [15:0] out_s119;
wire  [15:0] out_s120;
wire  [15:0] out_s121;
wire  [15:0] out_s122;
wire  [15:0] out_s123;
wire  [15:0] out_s124;
wire  [15:0] out_s125;
wire  [15:0] out_s126;
wire  [15:0] out_s127;
wire  [15:0] out_s128;
wire  [15:0] out_s129;
wire  [15:0] out_s130;
wire  [15:0] out_s131;
wire  [15:0] out_s132;
wire  [15:0] out_s133;
wire  [15:0] out_s134;
wire  [15:0] out_s135;
wire  [15:0] out_s136;
wire  [15:0] out_s137;
wire  [15:0] out_s138;
wire  [15:0] out_s139;
wire  [15:0] out_s140;
wire  [15:0] out_s141;
wire  [15:0] out_s142;
wire  [15:0] out_s143;
wire  [15:0] out_s144;
wire  [15:0] out_s145;
wire  [15:0] out_s146;
wire  [15:0] out_s147;
wire  [15:0] out_s148;
wire  [15:0] out_s149;
wire  [15:0] out_s150;
wire  [15:0] out_s151;
wire  [15:0] out_s152;
wire  [15:0] out_s153;
wire  [15:0] out_s154;
wire  [15:0] out_s155;
wire  [15:0] out_s156;
wire  [15:0] out_s157;
wire  [15:0] out_s158;
wire  [15:0] out_s159;
wire  [15:0] out_s160;
wire  [15:0] out_s161;
wire  [15:0] out_s162;
wire  [15:0] out_s163;
wire  [15:0] out_s164;
wire  [15:0] out_s165;
wire  [15:0] out_s166;
wire  [15:0] out_s167;
wire  [15:0] out_s168;
wire  [15:0] out_s169;
wire  [15:0] out_s170;
wire  [15:0] out_s171;
wire  [15:0] out_s172;
wire  [15:0] out_s173;
wire  [15:0] out_s174;
wire  [15:0] out_s175;
wire  [15:0] out_s176;
wire  [15:0] out_s177;
wire  [15:0] out_s178;
wire  [15:0] out_s179;
wire  [15:0] out_s180;
wire  [15:0] out_s181;
wire  [15:0] out_s182;
wire  [15:0] out_s183;
wire  [15:0] out_s184;
wire  [15:0] out_s185;
wire  [15:0] out_s186;
wire  [15:0] out_s187;
wire  [15:0] out_s188;
wire  [15:0] out_s189;
wire  [15:0] out_s190;
wire  [15:0] out_s191;
wire  [15:0] out_s192;
wire  [15:0] out_s193;
wire  [15:0] out_s194;
wire  [15:0] out_s195;
wire  [15:0] out_s196;
wire  [15:0] out_s197;
wire  [15:0] out_s198;
wire  [15:0] out_s199;
wire  [15:0] out_s200;
wire  [15:0] out_s201;
wire  [15:0] out_s202;
wire  [15:0] out_s203;
wire  [15:0] out_s204;
wire  [15:0] out_s205;
wire  [15:0] out_s206;
wire  [15:0] out_s207;
wire  [15:0] out_s208;
wire  [15:0] out_s209;
wire  [15:0] out_s210;
wire  [15:0] out_s211;
wire  [15:0] out_s212;
wire  [15:0] out_s213;
wire  [15:0] out_s214;
wire  [15:0] out_s215;
wire  [15:0] out_s216;
wire  [15:0] out_s217;
wire  [15:0] out_s218;
wire  [15:0] out_s219;
wire  [15:0] out_s220;
wire  [15:0] out_s221;
wire  [15:0] out_s222;
wire  [15:0] out_s223;
wire  [15:0] out_s224;
wire  [15:0] out_s225;
wire  [15:0] out_s226;
wire  [15:0] out_s227;
wire  [15:0] out_s228;
wire  [15:0] out_s229;
wire  [15:0] out_s230;
wire  [15:0] out_s231;
wire  [15:0] out_s232;
wire  [15:0] out_s233;
wire  [15:0] out_s234;
wire  [15:0] out_s235;
wire  [15:0] out_s236;
wire  [15:0] out_s237;
wire  [15:0] out_s238;
wire  [15:0] out_s239;
wire  [15:0] out_s240;
wire  [15:0] out_s241;
wire  [15:0] out_s242;
wire  [15:0] out_s243;
wire  [15:0] out_s244;
wire  [15:0] out_s245;
wire  [15:0] out_s246;
wire  [15:0] out_s247;
wire  [15:0] out_s248;
wire  [15:0] out_s249;
wire  [15:0] out_s250;
wire  [15:0] out_s251;
wire  [15:0] out_s252;
wire  [15:0] out_s253;
wire  [15:0] out_s254;
wire  [15:0] out_s255;
wire  [15:0] out_s256;
wire  [15:0] out_s257;
wire  [15:0] out_s258;
wire  [15:0] out_s259;
wire  [15:0] out_s260;
wire  [15:0] out_s261;
wire  [15:0] out_s262;
wire  [15:0] out_s263;
wire  [15:0] out_s264;
wire  [15:0] out_s265;
wire  [15:0] out_s266;
wire  [15:0] out_s267;
wire  [15:0] out_s268;
wire  [15:0] out_s269;
wire  [15:0] out_s270;
wire  [15:0] out_s271;
wire  [15:0] out_s272;
wire  [15:0] out_s273;
wire  [15:0] out_s274;
wire  [15:0] out_s275;
wire  [15:0] out_s276;
wire  [15:0] out_s277;
wire  [15:0] out_s278;
wire  [15:0] out_s279;
wire  [15:0] out_s280;
wire  [15:0] out_s281;
wire  [15:0] out_s282;
wire  [15:0] out_s283;
wire  [15:0] out_s284;
wire  [15:0] out_s285;
wire  [15:0] out_s286;
wire  [15:0] out_s287;
wire  [15:0] out_s288;
wire  [15:0] out_s289;
wire  [15:0] out_s290;
wire  [15:0] out_s291;
wire  [15:0] out_s292;
wire  [15:0] out_s293;
wire  [15:0] out_s294;
wire  [15:0] out_s295;
wire  [15:0] out_s296;
wire  [15:0] out_s297;
wire  [15:0] out_s298;
wire  [15:0] out_s299;
wire  [15:0] out_s300;
wire  [15:0] out_s301;
wire  [15:0] out_s302;
wire  [15:0] out_s303;
wire  [15:0] out_s304;
wire  [15:0] out_s305;
wire  [15:0] out_s306;
wire  [15:0] out_s307;
wire  [15:0] out_s308;
wire  [15:0] out_s309;
wire  [15:0] out_s310;
wire  [15:0] out_s311;
wire  [15:0] out_s312;
wire  [15:0] out_s313;
wire  [15:0] out_s314;
wire  [15:0] out_s315;
wire  [15:0] out_s316;
wire  [15:0] out_s317;
wire  [15:0] out_s318;
wire  [15:0] out_s319;
wire  [15:0] out_s320;
wire  [15:0] out_s321;
wire  [15:0] out_s322;
wire  [15:0] out_s323;
wire  [15:0] out_s324;
wire  [15:0] out_s325;
wire  [15:0] out_s326;
wire  [15:0] out_s327;
wire  [15:0] out_s328;
wire  [15:0] out_s329;
wire  [15:0] out_s330;
wire  [15:0] out_s331;
wire  [15:0] out_s332;
wire  [15:0] out_s333;
wire  [15:0] out_s334;
wire  [15:0] out_s335;
wire  [15:0] out_s336;
wire  [15:0] out_s337;
wire  [15:0] out_s338;
wire  [15:0] out_s339;
wire  [15:0] out_s340;
wire  [15:0] out_s341;
wire  [15:0] out_s342;
wire  [15:0] out_s343;
wire  [15:0] out_s344;
wire  [15:0] out_s345;
wire  [15:0] out_s346;
wire  [15:0] out_s347;
wire  [15:0] out_s348;
wire  [15:0] out_s349;
wire  [15:0] out_s350;
wire  [15:0] out_s351;
wire  [15:0] out_s352;
wire  [15:0] out_s353;
wire  [15:0] out_s354;
wire  [15:0] out_s355;
wire  [15:0] out_s356;
wire  [15:0] out_s357;
wire  [15:0] out_s358;
wire  [15:0] out_s359;
wire  [15:0] out_s360;
wire  [15:0] out_s361;
wire  [15:0] out_s362;
wire  [15:0] out_s363;
wire  [15:0] out_s364;
wire  [15:0] out_s365;
wire  [15:0] out_s366;
wire  [15:0] out_s367;
wire  [15:0] out_s368;
wire  [15:0] out_s369;
wire  [15:0] out_s370;
wire  [15:0] out_s371;
wire  [15:0] out_s372;
wire  [15:0] out_s373;
wire  [15:0] out_s374;
wire  [15:0] out_s375;
wire  [15:0] out_s376;
wire  [15:0] out_s377;
wire  [15:0] out_s378;
wire  [15:0] out_s379;
wire  [15:0] out_s380;
wire  [15:0] out_s381;
wire  [15:0] out_s382;
wire  [15:0] out_s383;
wire  [15:0] out_s384;
wire  [15:0] out_s385;
wire  [15:0] out_s386;
wire  [15:0] out_s387;
wire  [15:0] out_s388;
wire  [15:0] out_s389;
wire  [15:0] out_s390;
wire  [15:0] out_s391;
wire  [15:0] out_s392;
wire  [15:0] out_s393;
wire  [15:0] out_s394;
wire  [15:0] out_s395;
wire  [15:0] out_s396;
wire  [15:0] out_s397;
wire  [15:0] out_s398;
wire  [15:0] out_s399;
wire  [15:0] out_s400;
wire  [15:0] out_s401;
wire  [15:0] out_s402;
wire  [15:0] out_s403;
wire  [15:0] out_s404;
wire  [15:0] out_s405;
wire  [15:0] out_s406;
wire  [15:0] out_s407;
wire  [15:0] out_s408;
wire  [15:0] out_s409;
wire  [15:0] out_s410;
wire  [15:0] out_s411;
wire  [15:0] out_s412;
wire  [15:0] out_s413;
wire  [15:0] out_s414;
wire  [15:0] out_s415;
wire  [15:0] out_s416;
wire  [15:0] out_s417;
wire  [15:0] out_s418;
wire  [15:0] out_s419;
wire  [15:0] out_s420;
wire  [15:0] out_s421;
wire  [15:0] out_s422;
wire  [15:0] out_s423;
wire  [15:0] out_s424;
wire  [15:0] out_s425;
wire  [15:0] out_s426;
wire  [15:0] out_s427;
wire  [15:0] out_s428;
wire  [15:0] out_s429;
wire  [15:0] out_s430;
wire  [15:0] out_s431;
wire  [15:0] out_s432;
wire  [15:0] out_s433;
wire  [15:0] out_s434;
wire  [15:0] out_s435;
wire  [15:0] out_s436;
wire  [15:0] out_s437;
wire  [15:0] out_s438;
wire  [15:0] out_s439;
wire  [15:0] out_s440;
wire  [15:0] out_s441;
wire  [15:0] out_s442;
wire  [15:0] out_s443;
wire  [15:0] out_s444;
wire  [15:0] out_s445;
wire  [15:0] out_s446;
wire  [15:0] out_s447;
wire  [15:0] out_s448;
wire  [15:0] out_s449;
wire  [15:0] out_s450;
wire  [15:0] out_s451;
wire  [15:0] out_s452;
wire  [15:0] out_s453;
wire  [15:0] out_s454;
wire  [15:0] out_s455;
wire  [15:0] out_s456;
wire  [15:0] out_s457;
wire  [15:0] out_s458;
wire  [15:0] out_s459;
wire  [15:0] out_s460;
wire  [15:0] out_s461;
wire  [15:0] out_s462;
wire  [15:0] out_s463;
wire  [15:0] out_s464;
wire  [15:0] out_s465;
wire  [15:0] out_s466;
wire  [15:0] out_s467;
wire  [15:0] out_s468;
wire  [15:0] out_s469;
wire  [15:0] out_s470;
wire  [15:0] out_s471;
wire  [15:0] out_s472;
wire  [15:0] out_s473;
wire  [15:0] out_s474;
wire  [15:0] out_s475;
wire  [15:0] out_s476;
wire  [15:0] out_s477;
wire  [15:0] out_s478;
wire  [15:0] out_s479;
wire  [15:0] out_s480;
wire  [15:0] out_s481;
wire  [15:0] out_s482;
wire  [15:0] out_s483;
wire  [15:0] out_s484;
wire  [15:0] out_s485;
wire  [15:0] out_s486;
wire  [15:0] out_s487;
wire  [15:0] out_s488;
wire  [15:0] out_s489;
wire  [15:0] out_s490;
wire  [15:0] out_s491;
wire  [15:0] out_s492;
wire  [15:0] out_s493;
wire  [15:0] out_s494;
wire  [15:0] out_s495;
wire  [15:0] out_s496;
wire  [15:0] out_s497;
wire  [15:0] out_s498;
wire  [15:0] out_s499;
wire  [15:0] out_s500;
wire  [15:0] out_s501;
wire  [15:0] out_s502;
wire  [15:0] out_s503;
wire  [15:0] out_s504;
wire  [15:0] out_s505;
wire  [15:0] out_s506;
wire  [15:0] out_s507;
wire  [15:0] out_s508;
wire  [15:0] out_s509;
wire  [15:0] out_s510;
wire  [15:0] out_s511;
wire  [15:0] out_s512;
wire  [15:0] out_s513;
wire  [15:0] out_s514;
wire  [15:0] out_s515;
wire  [15:0] out_s516;
wire  [15:0] out_s517;
wire  [15:0] out_s518;
wire  [15:0] out_s519;
wire  [15:0] out_s520;
wire  [15:0] out_s521;
wire  [15:0] out_s522;
wire  [15:0] out_s523;
wire  [15:0] out_s524;
wire  [15:0] out_s525;
wire  [15:0] out_s526;
wire  [15:0] out_s527;
wire  [15:0] out_s528;
wire  [15:0] out_s529;
wire  [15:0] out_s530;
wire  [15:0] out_s531;
wire  [15:0] out_s532;
wire  [15:0] out_s533;
wire  [15:0] out_s534;
wire  [15:0] out_s535;
wire  [15:0] out_s536;
wire  [15:0] out_s537;
wire  [15:0] out_s538;
wire  [15:0] out_s539;
wire  [15:0] out_s540;
wire  [15:0] out_s541;
wire  [15:0] out_s542;
wire  [15:0] out_s543;
wire  [15:0] out_s544;
wire  [15:0] out_s545;
wire  [15:0] out_s546;
wire  [15:0] out_s547;
wire  [15:0] out_s548;
wire  [15:0] out_s549;
wire  [15:0] out_s550;
wire  [15:0] out_s551;
wire  [15:0] out_s552;
wire  [15:0] out_s553;
wire  [15:0] out_s554;
wire  [15:0] out_s555;
wire  [15:0] out_s556;
wire  [15:0] out_s557;
wire  [15:0] out_s558;
wire  [15:0] out_s559;
wire  [15:0] out_s560;
wire  [15:0] out_s561;
wire  [15:0] out_s562;
wire  [15:0] out_s563;
wire  [15:0] out_s564;
wire  [15:0] out_s565;
wire  [15:0] out_s566;
wire  [15:0] out_s567;
wire  [15:0] out_s568;
wire  [15:0] out_s569;
wire  [15:0] out_s570;
wire  [15:0] out_s571;
wire  [15:0] out_s572;
wire  [15:0] out_s573;
wire  [15:0] out_s574;
wire  [15:0] out_s575;
wire  [15:0] out_s576;
wire  [15:0] out_s577;
wire  [15:0] out_s578;
wire  [15:0] out_s579;
wire  [15:0] out_s580;
wire  [15:0] out_s581;
wire  [15:0] out_s582;
wire  [15:0] out_s583;
wire  [15:0] out_s584;
wire  [15:0] out_s585;
wire  [15:0] out_s586;
wire  [15:0] out_s587;
wire  [15:0] out_s588;
wire  [15:0] out_s589;
wire  [15:0] out_s590;
wire  [15:0] out_s591;
wire  [15:0] out_s592;
wire  [15:0] out_s593;
wire  [15:0] out_s594;
wire  [15:0] out_s595;
wire  [15:0] out_s596;
wire  [15:0] out_s597;
wire  [15:0] out_s598;
wire  [15:0] out_s599;
wire  [15:0] out_s600;
wire  [15:0] out_s601;
wire  [15:0] out_s602;
wire  [15:0] out_s603;
wire  [15:0] out_s604;
wire  [15:0] out_s605;
wire  [15:0] out_s606;
wire  [15:0] out_s607;
wire  [15:0] out_s608;
wire  [15:0] out_s609;
wire  [15:0] out_s610;
wire  [15:0] out_s611;
wire  [15:0] out_s612;
wire  [15:0] out_s613;
wire  [15:0] out_s614;
wire  [15:0] out_s615;
wire  [15:0] out_s616;
wire  [15:0] out_s617;
wire  [15:0] out_s618;
wire  [15:0] out_s619;
wire  [15:0] out_s620;
wire  [15:0] out_s621;
wire  [15:0] out_s622;
wire  [15:0] out_s623;
wire  [15:0] out_s624;
wire  [15:0] out_s625;
wire  [15:0] out_s626;
wire  [15:0] out_s627;
wire  [15:0] out_s628;
wire  [15:0] out_s629;
wire  [15:0] out_s630;
wire  [15:0] out_s631;
wire  [15:0] out_s632;
wire  [15:0] out_s633;
wire  [15:0] out_s634;
wire  [15:0] out_s635;
wire  [15:0] out_s636;
wire  [15:0] out_s637;
wire  [15:0] out_s638;
wire  [15:0] out_s639;
wire  [15:0] out_s640;
wire  [15:0] out_s641;
wire  [15:0] out_s642;
wire  [15:0] out_s643;
wire  [15:0] out_s644;
wire  [15:0] out_s645;
wire  [15:0] out_s646;
wire  [15:0] out_s647;
wire  [15:0] out_s648;
wire  [15:0] out_s649;
wire  [15:0] out_s650;
wire  [15:0] out_s651;
wire  [15:0] out_s652;
wire  [15:0] out_s653;
wire  [15:0] out_s654;
wire  [15:0] out_s655;
wire  [15:0] out_s656;
wire  [15:0] out_s657;
wire  [15:0] out_s658;
wire  [15:0] out_s659;
wire  [15:0] out_s660;
wire  [15:0] out_s661;
wire  [15:0] out_s662;
wire  [15:0] out_s663;
wire  [15:0] out_s664;
wire  [15:0] out_s665;
wire  [15:0] out_s666;
wire  [15:0] out_s667;
wire  [15:0] out_s668;
wire  [15:0] out_s669;
wire  [15:0] out_s670;
wire  [15:0] out_s671;
wire  [15:0] out_s672;
wire  [15:0] out_s673;
wire  [15:0] out_s674;
wire  [15:0] out_s675;
wire  [15:0] out_s676;
wire  [15:0] out_s677;
wire  [15:0] out_s678;
wire  [15:0] out_s679;
wire  [15:0] out_s680;
wire  [15:0] out_s681;
wire  [15:0] out_s682;
wire  [15:0] out_s683;
wire  [15:0] out_s684;
wire  [15:0] out_s685;
wire  [15:0] out_s686;
wire  [15:0] out_s687;
wire  [15:0] out_s688;
wire  [15:0] out_s689;
wire  [15:0] out_s690;
wire  [15:0] out_s691;
wire  [15:0] out_s692;
wire  [15:0] out_s693;
wire  [15:0] out_s694;
wire  [15:0] out_s695;
wire  [15:0] out_s696;
wire  [15:0] out_s697;
wire  [15:0] out_s698;
wire  [15:0] out_s699;
wire  [15:0] out_s700;
wire  [15:0] out_s701;
wire  [15:0] out_s702;
wire  [15:0] out_s703;
wire  [15:0] out_s704;
wire  [15:0] out_s705;
wire  [15:0] out_s706;
wire  [15:0] out_s707;
wire  [15:0] out_s708;
wire  [15:0] out_s709;
wire  [15:0] out_s710;
wire  [15:0] out_s711;
wire  [15:0] out_s712;
wire  [15:0] out_s713;
wire  [15:0] out_s714;
wire  [15:0] out_s715;
wire  [15:0] out_s716;
wire  [15:0] out_s717;
wire  [15:0] out_s718;
wire  [15:0] out_s719;
wire  [15:0] out_s720;
wire  [15:0] out_s721;
wire  [15:0] out_s722;
wire  [15:0] out_s723;
wire  [15:0] out_s724;
wire  [15:0] out_s725;
wire  [15:0] out_s726;
wire  [15:0] out_s727;
wire  [15:0] out_s728;
wire  [15:0] out_s729;
wire  [15:0] out_s730;
wire  [15:0] out_s731;
wire  [15:0] out_s732;
wire  [15:0] out_s733;
wire  [15:0] out_s734;
wire  [15:0] out_s735;
wire  [15:0] out_s736;
wire  [15:0] out_s737;
wire  [15:0] out_s738;
wire  [15:0] out_s739;
wire  [15:0] out_s740;
wire  [15:0] out_s741;
wire  [15:0] out_s742;
wire  [15:0] out_s743;
wire  [15:0] out_s744;
wire  [15:0] out_s745;
wire  [15:0] out_s746;
wire  [15:0] out_s747;
wire  [15:0] out_s748;
wire  [15:0] out_s749;
wire  [15:0] out_s750;
wire  [15:0] out_s751;
wire  [15:0] out_s752;
wire  [15:0] out_s753;
wire  [15:0] out_s754;
wire  [15:0] out_s755;
wire  [15:0] out_s756;
wire  [15:0] out_s757;
wire  [15:0] out_s758;
wire  [15:0] out_s759;
wire  [15:0] out_s760;
wire  [15:0] out_s761;
wire  [15:0] out_s762;
wire  [15:0] out_s763;
wire  [15:0] out_s764;
wire  [15:0] out_s765;
wire  [15:0] out_s766;
wire  [15:0] out_s767;
wire  [15:0] out_s768;
wire  [15:0] out_s769;
wire  [15:0] out_s770;
wire  [15:0] out_s771;
wire  [15:0] out_s772;
wire  [15:0] out_s773;
wire  [15:0] out_s774;
wire  [15:0] out_s775;
wire  [15:0] out_s776;
wire  [15:0] out_s777;
wire  [15:0] out_s778;
wire  [15:0] out_s779;
wire  [15:0] out_s780;
wire  [15:0] out_s781;
wire  [15:0] out_s782;
wire  [15:0] out_s783;
wire  [15:0] out_s784;
wire  [15:0] out_s785;
wire  [15:0] out_s786;
wire  [15:0] out_s787;
wire  [15:0] out_s788;
wire  [15:0] out_s789;
wire  [15:0] out_s790;
wire  [15:0] out_s791;
wire  [15:0] out_s792;
wire  [15:0] out_s793;
wire  [15:0] out_s794;
wire  [15:0] out_s795;
wire  [15:0] out_s796;
wire  [15:0] out_s797;
wire  [15:0] out_s798;
wire  [15:0] out_s799;
wire  [15:0] out_s800;
wire  [15:0] out_s801;
wire  [15:0] out_s802;
wire  [15:0] out_s803;
wire  [15:0] out_s804;
wire  [15:0] out_s805;
wire  [15:0] out_s806;
wire  [15:0] out_s807;
wire  [15:0] out_s808;
wire  [15:0] out_s809;
wire  [15:0] out_s810;
wire  [15:0] out_s811;
wire  [15:0] out_s812;
wire  [15:0] out_s813;
wire  [15:0] out_s814;
wire  [15:0] out_s815;
wire  [15:0] out_s816;
wire  [15:0] out_s817;
wire  [15:0] out_s818;
wire  [15:0] out_s819;
wire  [15:0] out_s820;
wire  [15:0] out_s821;
wire  [15:0] out_s822;
wire  [15:0] out_s823;
wire  [15:0] out_s824;
wire  [15:0] out_s825;
wire  [15:0] out_s826;
wire  [15:0] out_s827;
wire  [15:0] out_s828;
wire  [15:0] out_s829;
wire  [15:0] out_s830;
wire  [15:0] out_s831;
wire  [15:0] out_s832;
wire  [15:0] out_s833;
wire  [15:0] out_s834;
wire  [15:0] out_s835;
wire  [15:0] out_s836;
wire  [15:0] out_s837;
wire  [15:0] out_s838;
wire  [15:0] out_s839;
wire  [15:0] out_s840;
wire  [15:0] out_s841;
wire  [15:0] out_s842;
wire  [15:0] out_s843;
wire  [15:0] out_s844;
wire  [15:0] out_s845;
wire  [15:0] out_s846;
wire  [15:0] out_s847;
wire  [15:0] out_s848;
wire  [15:0] out_s849;
wire  [15:0] out_s850;
wire  [15:0] out_s851;
wire  [15:0] out_s852;
wire  [15:0] out_s853;
wire  [15:0] out_s854;
wire  [15:0] out_s855;
wire  [15:0] out_s856;
wire  [15:0] out_s857;
wire  [15:0] out_s858;
wire  [15:0] out_s859;
wire  [15:0] out_s860;
wire  [15:0] out_s861;
wire  [15:0] out_s862;
wire  [15:0] out_s863;
wire  [15:0] out_s864;
wire  [15:0] out_s865;
wire  [15:0] out_s866;
wire  [15:0] out_s867;
wire  [15:0] out_s868;
wire  [15:0] out_s869;
wire  [15:0] out_s870;
wire  [15:0] out_s871;
wire  [15:0] out_s872;
wire  [15:0] out_s873;
wire  [15:0] out_s874;
wire  [15:0] out_s875;
wire  [15:0] out_s876;
wire  [15:0] out_s877;
wire  [15:0] out_s878;
wire  [15:0] out_s879;
wire  [15:0] out_s880;
wire  [15:0] out_s881;
wire  [15:0] out_s882;
wire  [15:0] out_s883;
wire  [15:0] out_s884;
wire  [15:0] out_s885;
wire  [15:0] out_s886;
wire  [15:0] out_s887;
wire  [15:0] out_s888;
wire  [15:0] out_s889;
wire  [15:0] out_s890;
wire  [15:0] out_s891;
wire  [15:0] out_s892;
wire  [15:0] out_s893;
wire  [15:0] out_s894;
wire  [15:0] out_s895;
wire  [15:0] out_s896;
wire  [15:0] out_s897;
wire  [15:0] out_s898;
wire  [15:0] out_s899;
wire  [15:0] out_s900;
wire  [15:0] out_s901;
wire  [15:0] out_s902;
wire  [15:0] out_s903;
wire  [15:0] out_s904;
wire  [15:0] out_s905;
wire  [15:0] out_s906;
wire  [15:0] out_s907;
wire  [15:0] out_s908;
wire  [15:0] out_s909;
wire  [15:0] out_s910;
wire  [15:0] out_s911;
wire  [15:0] out_s912;
wire  [15:0] out_s913;
wire  [15:0] out_s914;
wire  [15:0] out_s915;
wire  [15:0] out_s916;
wire  [15:0] out_s917;
wire  [15:0] out_s918;
wire  [15:0] out_s919;
wire  [15:0] out_s920;
wire  [15:0] out_s921;
wire  [15:0] out_s922;
wire  [15:0] out_s923;
wire  [15:0] out_s924;
wire  [15:0] out_s925;
wire  [15:0] out_s926;
wire  [15:0] out_s927;
wire  [15:0] out_s928;
wire  [15:0] out_s929;
wire  [15:0] out_s930;
wire  [15:0] out_s931;
wire  [15:0] out_s932;
wire  [15:0] out_s933;
wire  [15:0] out_s934;
wire  [15:0] out_s935;
wire  [15:0] out_s936;
wire  [15:0] out_s937;
wire  [15:0] out_s938;
wire  [15:0] out_s939;
wire  [15:0] out_s940;
wire  [15:0] out_s941;
wire  [15:0] out_s942;
wire  [15:0] out_s943;
wire  [15:0] out_s944;
wire  [15:0] out_s945;
wire  [15:0] out_s946;
wire  [15:0] out_s947;
wire  [15:0] out_s948;
wire  [15:0] out_s949;
wire  [15:0] out_s950;
wire  [15:0] out_s951;
wire  [15:0] out_s952;
wire  [15:0] out_s953;
wire  [15:0] out_s954;
wire  [15:0] out_s955;
wire  [15:0] out_s956;
wire  [15:0] out_s957;
wire  [15:0] out_s958;
wire  [15:0] out_s959;
wire  [15:0] out_s960;
wire  [15:0] out_s961;
wire  [15:0] out_s962;
wire  [15:0] out_s963;
wire  [15:0] out_s964;
wire  [15:0] out_s965;
wire  [15:0] out_s966;
wire  [15:0] out_s967;
wire  [15:0] out_s968;
wire  [15:0] out_s969;
wire  [15:0] out_s970;
wire  [15:0] out_s971;
wire  [15:0] out_s972;
wire  [15:0] out_s973;
wire  [15:0] out_s974;
wire  [15:0] out_s975;
wire  [15:0] out_s976;
wire  [15:0] out_s977;
wire  [15:0] out_s978;
wire  [15:0] out_s979;
wire  [15:0] out_s980;
wire  [15:0] out_s981;
wire  [15:0] out_s982;
wire  [15:0] out_s983;
wire  [15:0] out_s984;
wire  [15:0] out_s985;
wire  [15:0] out_s986;
wire  [15:0] out_s987;
wire  [15:0] out_s988;
wire  [15:0] out_s989;
wire  [15:0] out_s990;
wire  [15:0] out_s991;
wire  [15:0] out_s992;
wire  [15:0] out_s993;
wire  [15:0] out_s994;
wire  [15:0] out_s995;
wire  [15:0] out_s996;
wire  [15:0] out_s997;
wire  [15:0] out_s998;
wire  [15:0] out_s999;
wire  [15:0] out_s1000;
wire  [15:0] out_s1001;
wire  [15:0] out_s1002;
wire  [15:0] out_s1003;
wire  [15:0] out_s1004;
wire  [15:0] out_s1005;
wire  [15:0] out_s1006;
wire  [15:0] out_s1007;
wire  [15:0] out_s1008;
wire  [15:0] out_s1009;
wire  [15:0] out_s1010;
wire  [15:0] out_s1011;
wire  [15:0] out_s1012;
wire  [15:0] out_s1013;
wire  [15:0] out_s1014;
wire  [15:0] out_s1015;
wire  [15:0] out_s1016;
wire  [15:0] out_s1017;
wire  [15:0] out_s1018;
wire  [15:0] out_s1019;
wire  [15:0] out_s1020;
wire  [15:0] out_s1021;
wire  [15:0] out_s1022;
wire  [15:0] out_s1023;
wire  [15:0] out_s1024;
wire  [15:0] out_s1025;
wire  [15:0] out_s1026;
wire  [15:0] out_s1027;
wire  [15:0] out_s1028;
wire  [15:0] out_s1029;
wire  [15:0] out_s1030;
wire  [15:0] out_s1031;
wire  [15:0] out_s1032;
wire  [15:0] out_s1033;
wire  [15:0] out_s1034;
wire  [15:0] out_s1035;
wire  [15:0] out_s1036;
wire  [15:0] out_s1037;
wire  [15:0] out_s1038;
wire  [15:0] out_s1039;
wire  [15:0] out_s1040;
wire  [15:0] out_s1041;
wire  [15:0] out_s1042;
wire  [15:0] out_s1043;
wire  [15:0] out_s1044;
wire  [15:0] out_s1045;
wire  [15:0] out_s1046;
wire  [15:0] out_s1047;
wire  [15:0] out_s1048;
wire  [15:0] out_s1049;
wire  [15:0] out_s1050;
wire  [15:0] out_s1051;
wire  [15:0] out_s1052;
wire  [15:0] out_s1053;
wire  [15:0] out_s1054;
wire  [15:0] out_s1055;
wire  [15:0] out_s1056;
wire  [15:0] out_s1057;
wire  [15:0] out_s1058;
wire  [15:0] out_s1059;
wire  [15:0] out_s1060;
wire  [15:0] out_s1061;
wire  [15:0] out_s1062;
wire  [15:0] out_s1063;
wire  [15:0] out_s1064;
wire  [15:0] out_s1065;
wire  [15:0] out_s1066;
wire  [15:0] out_s1067;
wire  [15:0] out_s1068;
wire  [15:0] out_s1069;
wire  [15:0] out_s1070;
wire  [15:0] out_s1071;
wire  [15:0] out_s1072;
wire  [15:0] out_s1073;
wire  [15:0] out_s1074;
wire  [15:0] out_s1075;
wire  [15:0] out_s1076;
wire  [15:0] out_s1077;
wire  [15:0] out_s1078;
wire  [15:0] out_s1079;
wire  [15:0] out_s1080;
wire  [15:0] out_s1081;
wire  [15:0] out_s1082;
wire  [15:0] out_s1083;
wire  [15:0] out_s1084;
wire  [15:0] out_s1085;
wire  [15:0] out_s1086;
wire  [15:0] out_s1087;
wire  [15:0] out_s1088;
wire  [15:0] out_s1089;
wire  [15:0] out_s1090;
wire  [15:0] out_s1091;
wire  [15:0] out_s1092;
wire  [15:0] out_s1093;
wire  [15:0] out_s1094;
wire  [15:0] out_s1095;
wire  [15:0] out_s1096;
wire  [15:0] out_s1097;
wire  [15:0] out_s1098;
wire  [15:0] out_s1099;
wire  [15:0] out_s1100;
wire  [15:0] out_s1101;
wire  [15:0] out_s1102;
wire  [15:0] out_s1103;
wire  [15:0] out_s1104;
wire  [15:0] out_s1105;
wire  [15:0] out_s1106;
wire  [15:0] out_s1107;
wire  [15:0] out_s1108;
wire  [15:0] out_s1109;
wire  [15:0] out_s1110;
wire  [15:0] out_s1111;
wire  [15:0] out_s1112;
wire  [15:0] out_s1113;
wire  [15:0] out_s1114;
wire  [15:0] out_s1115;
wire  [15:0] out_s1116;
wire  [15:0] out_s1117;
wire  [15:0] out_s1118;
wire  [15:0] out_s1119;
wire  [15:0] out_s1120;
wire  [15:0] out_s1121;
wire  [15:0] out_s1122;
wire  [15:0] out_s1123;
wire  [15:0] out_s1124;
wire  [15:0] out_s1125;
wire  [15:0] out_s1126;
wire  [15:0] out_s1127;
wire  [15:0] out_s1128;
wire  [15:0] out_s1129;
wire  [15:0] out_s1130;
wire  [15:0] out_s1131;
wire  [15:0] out_s1132;
wire  [15:0] out_s1133;
wire  [15:0] out_s1134;
wire  [15:0] out_s1135;
wire  [15:0] out_s1136;
wire  [15:0] out_s1137;
wire  [15:0] out_s1138;
wire  [15:0] out_s1139;
wire  [15:0] out_s1140;
wire  [15:0] out_s1141;
wire  [15:0] out_s1142;
wire  [15:0] out_s1143;
wire  [15:0] out_s1144;
wire  [15:0] out_s1145;
wire  [15:0] out_s1146;
wire  [15:0] out_s1147;
wire  [15:0] out_s1148;
wire  [15:0] out_s1149;
wire  [15:0] out_s1150;
wire  [15:0] out_s1151;
wire  [15:0] out_s1152;
wire  [15:0] out_s1153;
wire  [15:0] out_s1154;
wire  [15:0] out_s1155;
wire  [15:0] out_s1156;
wire  [15:0] out_s1157;
wire  [15:0] out_s1158;
wire  [15:0] out_s1159;
wire  [15:0] out_s1160;
wire  [15:0] out_s1161;
wire  [15:0] out_s1162;
wire  [15:0] out_s1163;
wire  [15:0] out_s1164;
wire  [15:0] out_s1165;
wire  [15:0] out_s1166;
wire  [15:0] out_s1167;
wire  [15:0] out_s1168;
wire  [15:0] out_s1169;
wire  [15:0] out_s1170;
wire  [15:0] out_s1171;
wire  [15:0] out_s1172;
wire  [15:0] out_s1173;
wire  [15:0] out_s1174;
wire  [15:0] out_s1175;
wire  [15:0] out_s1176;
wire  [15:0] out_s1177;
wire  [15:0] out_s1178;
wire  [15:0] out_s1179;
wire  [15:0] out_s1180;
wire  [15:0] out_s1181;
wire  [15:0] out_s1182;
wire  [15:0] out_s1183;
wire  [15:0] out_s1184;
wire  [15:0] out_s1185;
wire  [15:0] out_s1186;
wire  [15:0] out_s1187;
wire  [15:0] out_s1188;
wire  [15:0] out_s1189;
wire  [15:0] out_s1190;
wire  [15:0] out_s1191;
wire  [15:0] out_s1192;
wire  [15:0] out_s1193;
wire  [15:0] out_s1194;
wire  [15:0] out_s1195;
wire  [15:0] out_s1196;
wire  [15:0] out_s1197;
wire  [15:0] out_s1198;
wire  [15:0] out_s1199;
wire  [15:0] out_s1200;
wire  [15:0] out_s1201;
wire  [15:0] out_s1202;
wire  [15:0] out_s1203;
wire  [15:0] out_s1204;
wire  [15:0] out_s1205;
wire  [15:0] out_s1206;
wire  [15:0] out_s1207;
wire  [15:0] out_s1208;
wire  [15:0] out_s1209;
wire  [15:0] out_s1210;
wire  [15:0] out_s1211;
wire  [15:0] out_s1212;
wire  [15:0] out_s1213;
wire  [15:0] out_s1214;
wire  [15:0] out_s1215;
wire  [15:0] out_s1216;
wire  [15:0] out_s1217;
wire  [15:0] out_s1218;
wire  [15:0] out_s1219;
wire  [15:0] out_s1220;
wire  [15:0] out_s1221;
wire  [15:0] out_s1222;
wire  [15:0] out_s1223;
wire  [15:0] out_s1224;
wire  [15:0] out_s1225;
wire  [15:0] out_s1226;
wire  [15:0] out_s1227;
wire  [15:0] out_s1228;
wire  [15:0] out_s1229;
wire  [15:0] out_s1230;
wire  [15:0] out_s1231;
wire  [15:0] out_s1232;
wire  [15:0] out_s1233;
wire  [15:0] out_s1234;
wire  [15:0] out_s1235;
wire  [15:0] out_s1236;
wire  [15:0] out_s1237;
wire  [15:0] out_s1238;
wire  [15:0] out_s1239;
wire  [15:0] out_s1240;
wire  [15:0] out_s1241;
wire  [15:0] out_s1242;
wire  [15:0] out_s1243;
wire  [15:0] out_s1244;
wire  [15:0] out_s1245;
wire  [15:0] out_s1246;
wire  [15:0] out_s1247;
wire  [15:0] out_s1248;
wire  [15:0] out_s1249;
wire  [15:0] out_s1250;
wire  [15:0] out_s1251;
wire  [15:0] out_s1252;
wire  [15:0] out_s1253;
wire  [15:0] out_s1254;
wire  [15:0] out_s1255;
wire  [15:0] out_s1256;
wire  [15:0] out_s1257;
wire  [15:0] out_s1258;
wire  [15:0] out_s1259;
wire  [15:0] out_s1260;
wire  [15:0] out_s1261;
wire  [15:0] out_s1262;
wire  [15:0] out_s1263;
wire  [15:0] out_s1264;
wire  [15:0] out_s1265;
wire  [15:0] out_s1266;
wire  [15:0] out_s1267;
wire  [15:0] out_s1268;
wire  [15:0] out_s1269;
wire  [15:0] out_s1270;
wire  [15:0] out_s1271;
wire  [15:0] out_s1272;
wire  [15:0] out_s1273;
wire  [15:0] out_s1274;
wire  [15:0] out_s1275;
wire  [15:0] out_s1276;
wire  [15:0] out_s1277;
wire  [15:0] out_s1278;
wire  [15:0] out_s1279;
wire  [15:0] out_s1280;
wire  [15:0] out_s1281;
wire  [15:0] out_s1282;
wire  [15:0] out_s1283;
wire  [15:0] out_s1284;
wire  [15:0] out_s1285;
wire  [15:0] out_s1286;
wire  [15:0] out_s1287;
wire  [15:0] out_s1288;
wire  [15:0] out_s1289;
wire  [15:0] out_s1290;
wire  [15:0] out_s1291;
wire  [15:0] out_s1292;
wire  [15:0] out_s1293;
wire  [15:0] out_s1294;
wire  [15:0] out_s1295;
wire  [15:0] out_s1296;
wire  [15:0] out_s1297;
wire  [15:0] out_s1298;
wire  [15:0] out_s1299;
wire  [15:0] out_s1300;
wire  [15:0] out_s1301;
wire  [15:0] out_s1302;
wire  [15:0] out_s1303;
wire  [15:0] out_s1304;
wire  [15:0] out_s1305;
wire  [15:0] out_s1306;
wire  [15:0] out_s1307;
wire  [15:0] out_s1308;
wire  [15:0] out_s1309;
wire  [15:0] out_s1310;
wire  [15:0] out_s1311;
wire  [15:0] out_s1312;
wire  [15:0] out_s1313;
wire  [15:0] out_s1314;
wire  [15:0] out_s1315;
wire  [15:0] out_s1316;
wire  [15:0] out_s1317;
wire  [15:0] out_s1318;
wire  [15:0] out_s1319;
wire  [15:0] out_s1320;
wire  [15:0] out_s1321;
wire  [15:0] out_s1322;
wire  [15:0] out_s1323;
wire  [15:0] out_s1324;
wire  [15:0] out_s1325;
wire  [15:0] out_s1326;
wire  [15:0] out_s1327;
wire  [15:0] out_s1328;
wire  [15:0] out_s1329;
wire  [15:0] out_s1330;
wire  [15:0] out_s1331;
wire  [15:0] out_s1332;
wire  [15:0] out_s1333;
wire  [15:0] out_s1334;
wire  [15:0] out_s1335;
wire  [15:0] out_s1336;
wire  [15:0] out_s1337;
wire  [15:0] out_s1338;
wire  [15:0] out_s1339;
wire  [15:0] out_s1340;
wire  [15:0] out_s1341;
wire  [15:0] out_s1342;
wire  [15:0] out_s1343;
wire  [15:0] out_s1344;
wire  [15:0] out_s1345;
wire  [15:0] out_s1346;
wire  [15:0] out_s1347;
wire  [15:0] out_s1348;
wire  [15:0] out_s1349;
wire  [15:0] out_s1350;
wire  [15:0] out_s1351;
wire  [15:0] out_s1352;
wire  [15:0] out_s1353;
wire  [15:0] out_s1354;
wire  [15:0] out_s1355;
wire  [15:0] out_s1356;
wire  [15:0] out_s1357;
wire  [15:0] out_s1358;
wire  [15:0] out_s1359;
wire  [15:0] out_s1360;
wire  [15:0] out_s1361;
wire  [15:0] out_s1362;
wire  [15:0] out_s1363;
wire  [15:0] out_s1364;
wire  [15:0] out_s1365;
wire  [15:0] out_s1366;
wire  [15:0] out_s1367;
wire  [15:0] out_s1368;
wire  [15:0] out_s1369;
wire  [15:0] out_s1370;
wire  [15:0] out_s1371;
wire  [15:0] out_s1372;
wire  [15:0] out_s1373;
wire  [15:0] out_s1374;
wire  [15:0] out_s1375;
wire  [15:0] out_s1376;
wire  [15:0] out_s1377;
wire  [15:0] out_s1378;
wire  [15:0] out_s1379;
wire  [15:0] out_s1380;
wire  [15:0] out_s1381;
wire  [15:0] out_s1382;
wire  [15:0] out_s1383;
wire  [15:0] out_s1384;
wire  [15:0] out_s1385;
wire  [15:0] out_s1386;
wire  [15:0] out_s1387;
wire  [15:0] out_s1388;
wire  [15:0] out_s1389;
wire  [15:0] out_s1390;
wire  [15:0] out_s1391;
wire  [15:0] out_s1392;
wire  [15:0] out_s1393;
wire  [15:0] out_s1394;
wire  [15:0] out_s1395;
wire  [15:0] out_s1396;
wire  [15:0] out_s1397;
wire  [15:0] out_s1398;
wire  [15:0] out_s1399;
wire  [15:0] out_s1400;
wire  [15:0] out_s1401;
wire  [15:0] out_s1402;
wire  [15:0] out_s1403;
wire  [15:0] out_s1404;
wire  [15:0] out_s1405;
wire  [15:0] out_s1406;
wire  [15:0] out_s1407;
wire  [15:0] out_s1408;
wire  [15:0] out_s1409;
wire  [15:0] out_s1410;
wire  [15:0] out_s1411;
wire  [15:0] out_s1412;
wire  [15:0] out_s1413;
wire  [15:0] out_s1414;
wire  [15:0] out_s1415;
wire  [15:0] out_s1416;
wire  [15:0] out_s1417;
wire  [15:0] out_s1418;
wire  [15:0] out_s1419;
wire  [15:0] out_s1420;
wire  [15:0] out_s1421;
wire  [15:0] out_s1422;
wire  [15:0] out_s1423;
wire  [15:0] out_s1424;
wire  [15:0] out_s1425;
wire  [15:0] out_s1426;
wire  [15:0] out_s1427;
wire  [15:0] out_s1428;
wire  [15:0] out_s1429;
wire  [15:0] out_s1430;
wire  [15:0] out_s1431;
wire  [15:0] out_s1432;
wire  [15:0] out_s1433;
wire  [15:0] out_s1434;
wire  [15:0] out_s1435;
wire  [15:0] out_s1436;
wire  [15:0] out_s1437;
wire  [15:0] out_s1438;
wire  [15:0] out_s1439;
wire  [15:0] out_s1440;
wire  [15:0] out_s1441;
wire  [15:0] out_s1442;
wire  [15:0] out_s1443;
wire  [15:0] out_s1444;
wire  [15:0] out_s1445;
wire  [15:0] out_s1446;
wire  [15:0] out_s1447;
wire  [15:0] out_s1448;
wire  [15:0] out_s1449;
wire  [15:0] out_s1450;
wire  [15:0] out_s1451;
wire  [15:0] out_s1452;
wire  [15:0] out_s1453;
wire  [15:0] out_s1454;
wire  [15:0] out_s1455;
wire  [15:0] out_s1456;
wire  [15:0] out_s1457;
wire  [15:0] out_s1458;
wire  [15:0] out_s1459;
wire  [15:0] out_s1460;
wire  [15:0] out_s1461;
wire  [15:0] out_s1462;
wire  [15:0] out_s1463;
wire  [15:0] out_s1464;
wire  [15:0] out_s1465;
wire  [15:0] out_s1466;
wire  [15:0] out_s1467;
wire  [15:0] out_s1468;
wire  [15:0] out_s1469;
wire  [15:0] out_s1470;
wire  [15:0] out_s1471;
wire  [15:0] out_s1472;
wire  [15:0] out_s1473;
wire  [15:0] out_s1474;
wire  [15:0] out_s1475;
wire  [15:0] out_s1476;
wire  [15:0] out_s1477;
wire  [15:0] out_s1478;
wire  [15:0] out_s1479;
wire  [15:0] out_s1480;
wire  [15:0] out_s1481;
wire  [15:0] out_s1482;
wire  [15:0] out_s1483;
wire  [15:0] out_s1484;
wire  [15:0] out_s1485;
wire  [15:0] out_s1486;
wire  [15:0] out_s1487;
wire  [15:0] out_s1488;
wire  [15:0] out_s1489;
wire  [15:0] out_s1490;
wire  [15:0] out_s1491;
wire  [15:0] out_s1492;
wire  [15:0] out_s1493;
wire  [15:0] out_s1494;
wire  [15:0] out_s1495;
wire  [15:0] out_s1496;
wire  [15:0] out_s1497;
wire  [15:0] out_s1498;
wire  [15:0] out_s1499;
wire  [15:0] out_s1500;
wire  [15:0] out_s1501;
wire  [15:0] out_s1502;
wire  [15:0] out_s1503;
wire  [15:0] out_s1504;
wire  [15:0] out_s1505;
wire  [15:0] out_s1506;
wire  [15:0] out_s1507;
wire  [15:0] out_s1508;
wire  [15:0] out_s1509;
wire  [15:0] out_s1510;
wire  [15:0] out_s1511;
wire  [15:0] out_s1512;
wire  [15:0] out_s1513;
wire  [15:0] out_s1514;
wire  [15:0] out_s1515;
wire  [15:0] out_s1516;
wire  [15:0] out_s1517;
wire  [15:0] out_s1518;
wire  [15:0] out_s1519;
wire  [15:0] out_s1520;
wire  [15:0] out_s1521;
wire  [15:0] out_s1522;
wire  [15:0] out_s1523;
wire  [15:0] out_s1524;
wire  [15:0] out_s1525;
wire  [15:0] out_s1526;
wire  [15:0] out_s1527;
wire  [15:0] out_s1528;
wire  [15:0] out_s1529;
wire  [15:0] out_s1530;
wire  [15:0] out_s1531;
wire  [15:0] out_s1532;
wire  [15:0] out_s1533;
wire  [15:0] out_s1534;
wire  [15:0] out_s1535;
wire  [15:0] out_s1536;
wire  [15:0] out_s1537;
wire  [15:0] out_s1538;
wire  [15:0] out_s1539;
wire  [15:0] out_s1540;
wire  [15:0] out_s1541;
wire  [15:0] out_s1542;
wire  [15:0] out_s1543;
wire  [15:0] out_s1544;
wire  [15:0] out_s1545;
wire  [15:0] out_s1546;
wire  [15:0] out_s1547;
wire  [15:0] out_s1548;
wire  [15:0] out_s1549;
wire  [15:0] out_s1550;
wire  [15:0] out_s1551;
wire  [15:0] out_s1552;
wire  [15:0] out_s1553;
wire  [15:0] out_s1554;
wire  [15:0] out_s1555;
wire  [15:0] out_s1556;
wire  [15:0] out_s1557;
wire  [15:0] out_s1558;
wire  [15:0] out_s1559;
wire  [15:0] out_s1560;
wire  [15:0] out_s1561;
wire  [15:0] out_s1562;
wire  [15:0] out_s1563;
wire  [15:0] out_s1564;
wire  [15:0] out_s1565;
wire  [15:0] out_s1566;
wire  [15:0] out_s1567;
wire  [15:0] out_s1568;
wire  [15:0] out_s1569;
wire  [15:0] out_s1570;
wire  [15:0] out_s1571;
wire  [15:0] out_s1572;
wire  [15:0] out_s1573;
wire  [15:0] out_s1574;
wire  [15:0] out_s1575;
wire  [15:0] out_s1576;
wire  [15:0] out_s1577;
wire  [15:0] out_s1578;
wire  [15:0] out_s1579;
wire  [15:0] out_s1580;
wire  [15:0] out_s1581;
wire  [15:0] out_s1582;
wire  [15:0] out_s1583;
wire  [15:0] out_s1584;
wire  [15:0] out_s1585;
wire  [15:0] out_s1586;
wire  [15:0] out_s1587;
wire  [15:0] out_s1588;
wire  [15:0] out_s1589;
wire  [15:0] out_s1590;
wire  [15:0] out_s1591;
wire  [15:0] out_s1592;
wire  [15:0] out_s1593;
wire  [15:0] out_s1594;
wire  [15:0] out_s1595;
wire  [15:0] out_s1596;
wire  [15:0] out_s1597;
wire  [15:0] out_s1598;
wire  [15:0] out_s1599;
wire  [15:0] out_s1600;
wire  [15:0] out_s1601;
wire  [15:0] out_s1602;
wire  [15:0] out_s1603;
wire  [15:0] out_s1604;
wire  [15:0] out_s1605;
wire  [15:0] out_s1606;
wire  [15:0] out_s1607;
wire  [15:0] out_s1608;
wire  [15:0] out_s1609;
wire  [15:0] out_s1610;
wire  [15:0] out_s1611;
wire  [15:0] out_s1612;
wire  [15:0] out_s1613;
wire  [15:0] out_s1614;
wire  [15:0] out_s1615;
wire  [15:0] out_s1616;
wire  [15:0] out_s1617;
wire  [15:0] out_s1618;
wire  [15:0] out_s1619;
wire  [15:0] out_s1620;
wire  [15:0] out_s1621;
wire  [15:0] out_s1622;
wire  [15:0] out_s1623;
wire  [15:0] out_s1624;
wire  [15:0] out_s1625;
wire  [15:0] out_s1626;
wire  [15:0] out_s1627;
wire  [15:0] out_s1628;
wire  [15:0] out_s1629;
wire  [15:0] out_s1630;
wire  [15:0] out_s1631;
wire  [15:0] out_s1632;
wire  [15:0] out_s1633;
wire  [15:0] out_s1634;
wire  [15:0] out_s1635;
wire  [15:0] out_s1636;
wire  [15:0] out_s1637;
wire  [15:0] out_s1638;
wire  [15:0] out_s1639;
wire  [15:0] out_s1640;
wire  [15:0] out_s1641;
wire  [15:0] out_s1642;
wire  [15:0] out_s1643;
wire  [15:0] out_s1644;
wire  [15:0] out_s1645;
wire  [15:0] out_s1646;
wire  [15:0] out_s1647;
wire  [15:0] out_s1648;
wire  [15:0] out_s1649;
wire  [15:0] out_s1650;
wire  [15:0] out_s1651;
wire  [15:0] out_s1652;
wire  [15:0] out_s1653;
wire  [15:0] out_s1654;
wire  [15:0] out_s1655;
wire  [15:0] out_s1656;
wire  [15:0] out_s1657;
wire  [15:0] out_s1658;
wire  [15:0] out_s1659;
wire  [15:0] out_s1660;
wire  [15:0] out_s1661;
wire  [15:0] out_s1662;
wire  [15:0] out_s1663;
wire  [15:0] out_s1664;
wire  [15:0] out_s1665;
wire  [15:0] out_s1666;
wire  [15:0] out_s1667;
wire  [15:0] out_s1668;
wire  [15:0] out_s1669;
wire  [15:0] out_s1670;
wire  [15:0] out_s1671;
wire  [15:0] out_s1672;
wire  [15:0] out_s1673;
wire  [15:0] out_s1674;
wire  [15:0] out_s1675;
wire  [15:0] out_s1676;
wire  [15:0] out_s1677;
wire  [15:0] out_s1678;
wire  [15:0] out_s1679;
wire  [15:0] out_s1680;
wire  [15:0] out_s1681;
wire  [15:0] out_s1682;
wire  [15:0] out_s1683;
wire  [15:0] out_s1684;
wire  [15:0] out_s1685;
wire  [15:0] out_s1686;
wire  [15:0] out_s1687;
wire  [15:0] out_s1688;
wire  [15:0] out_s1689;
wire  [15:0] out_s1690;
wire  [15:0] out_s1691;
wire  [15:0] out_s1692;
wire  [15:0] out_s1693;
wire  [15:0] out_s1694;
wire  [15:0] out_s1695;
wire  [15:0] out_s1696;
wire  [15:0] out_s1697;
wire  [15:0] out_s1698;
wire  [15:0] out_s1699;
wire  [15:0] out_s1700;
wire  [15:0] out_s1701;
wire  [15:0] out_s1702;
wire  [15:0] out_s1703;
wire  [15:0] out_s1704;
wire  [15:0] out_s1705;
wire  [15:0] out_s1706;
wire  [15:0] out_s1707;
wire  [15:0] out_s1708;
wire  [15:0] out_s1709;
wire  [15:0] out_s1710;
wire  [15:0] out_s1711;
wire  [15:0] out_s1712;
wire  [15:0] out_s1713;
wire  [15:0] out_s1714;
wire  [15:0] out_s1715;
wire  [15:0] out_s1716;
wire  [15:0] out_s1717;
wire  [15:0] out_s1718;
wire  [15:0] out_s1719;
wire  [15:0] out_s1720;
wire  [15:0] out_s1721;
wire  [15:0] out_s1722;
wire  [15:0] out_s1723;
wire  [15:0] out_s1724;
wire  [15:0] out_s1725;
wire  [15:0] out_s1726;
wire  [15:0] out_s1727;
wire  [15:0] out_s1728;
wire  [15:0] out_s1729;
wire  [15:0] out_s1730;
wire  [15:0] out_s1731;
wire  [15:0] out_s1732;
wire  [15:0] out_s1733;
wire  [15:0] out_s1734;
wire  [15:0] out_s1735;
wire  [15:0] out_s1736;
wire  [15:0] out_s1737;
wire  [15:0] out_s1738;
wire  [15:0] out_s1739;
wire  [15:0] out_s1740;
wire  [15:0] out_s1741;
wire  [15:0] out_s1742;
wire  [15:0] out_s1743;
wire  [15:0] out_s1744;
wire  [15:0] out_s1745;
wire  [15:0] out_s1746;
wire  [15:0] out_s1747;
wire  [15:0] out_s1748;
wire  [15:0] out_s1749;
wire  [15:0] out_s1750;
wire  [15:0] out_s1751;
wire  [15:0] out_s1752;
wire  [15:0] out_s1753;
wire  [15:0] out_s1754;
wire  [15:0] out_s1755;
wire  [15:0] out_s1756;
wire  [15:0] out_s1757;
wire  [15:0] out_s1758;
wire  [15:0] out_s1759;
wire  [15:0] out_s1760;
wire  [15:0] out_s1761;
wire  [15:0] out_s1762;
wire  [15:0] out_s1763;
wire  [15:0] out_s1764;
wire  [15:0] out_s1765;
wire  [15:0] out_s1766;
wire  [15:0] out_s1767;
wire  [15:0] out_s1768;
wire  [15:0] out_s1769;
wire  [15:0] out_s1770;
wire  [15:0] out_s1771;
wire  [15:0] out_s1772;
wire  [15:0] out_s1773;
wire  [15:0] out_s1774;
wire  [15:0] out_s1775;
wire  [15:0] out_s1776;
wire  [15:0] out_s1777;
wire  [15:0] out_s1778;
wire  [15:0] out_s1779;
wire  [15:0] out_s1780;
wire  [15:0] out_s1781;
wire  [15:0] out_s1782;
wire  [15:0] out_s1783;
wire  [15:0] out_s1784;
wire  [15:0] out_s1785;
wire  [15:0] out_s1786;
wire  [15:0] out_s1787;
wire  [15:0] out_s1788;
wire  [15:0] out_s1789;
wire  [15:0] out_s1790;
wire  [15:0] out_s1791;
wire  [15:0] out_s1792;
wire  [15:0] out_s1793;
wire  [15:0] out_s1794;
wire  [15:0] out_s1795;
wire  [15:0] out_s1796;
wire  [15:0] out_s1797;
wire  [15:0] out_s1798;
wire  [15:0] out_s1799;
wire  [15:0] out_s1800;
wire  [15:0] out_s1801;
wire  [15:0] out_s1802;
wire  [15:0] out_s1803;
wire  [15:0] out_s1804;
wire  [15:0] out_s1805;
wire  [15:0] out_s1806;
wire  [15:0] out_s1807;
wire  [15:0] out_s1808;
wire  [15:0] out_s1809;
wire  [15:0] out_s1810;
wire  [15:0] out_s1811;
wire  [15:0] out_s1812;
wire  [15:0] out_s1813;
wire  [15:0] out_s1814;
wire  [15:0] out_s1815;
wire  [15:0] out_s1816;
wire  [15:0] out_s1817;
wire  [15:0] out_s1818;
wire  [15:0] out_s1819;
wire  [15:0] out_s1820;
wire  [15:0] out_s1821;
wire  [15:0] out_s1822;
wire  [15:0] out_s1823;
wire  [15:0] out_s1824;
wire  [15:0] out_s1825;
wire  [15:0] out_s1826;
wire  [15:0] out_s1827;
wire  [15:0] out_s1828;
wire  [15:0] out_s1829;
wire  [15:0] out_s1830;
wire  [15:0] out_s1831;
wire  [15:0] out_s1832;
wire  [15:0] out_s1833;
wire  [15:0] out_s1834;
wire  [15:0] out_s1835;
wire  [15:0] out_s1836;
wire  [15:0] out_s1837;
wire  [15:0] out_s1838;
wire  [15:0] out_s1839;
wire  [15:0] out_s1840;
wire  [15:0] out_s1841;
wire  [15:0] out_s1842;
wire  [15:0] out_s1843;
wire  [15:0] out_s1844;
wire  [15:0] out_s1845;
wire  [15:0] out_s1846;
wire  [15:0] out_s1847;
wire  [15:0] out_s1848;
wire  [15:0] out_s1849;
wire  [15:0] out_s1850;
wire  [15:0] out_s1851;
wire  [15:0] out_s1852;
wire  [15:0] out_s1853;
wire  [15:0] out_s1854;
wire  [15:0] out_s1855;
wire  [15:0] out_s1856;
wire  [15:0] out_s1857;
wire  [15:0] out_s1858;
wire  [15:0] out_s1859;
wire  [15:0] out_s1860;
wire  [15:0] out_s1861;
wire  [15:0] out_s1862;
wire  [15:0] out_s1863;
wire  [15:0] out_s1864;
wire  [15:0] out_s1865;
wire  [15:0] out_s1866;
wire  [15:0] out_s1867;
wire  [15:0] out_s1868;
wire  [15:0] out_s1869;
wire  [15:0] out_s1870;
wire  [15:0] out_s1871;
wire  [15:0] out_s1872;
wire  [15:0] out_s1873;
wire  [15:0] out_s1874;
wire  [15:0] out_s1875;
wire  [15:0] out_s1876;
wire  [15:0] out_s1877;
wire  [15:0] out_s1878;
wire  [15:0] out_s1879;
wire  [15:0] out_s1880;
wire  [15:0] out_s1881;
wire  [15:0] out_s1882;
wire  [15:0] out_s1883;
wire  [15:0] out_s1884;
wire  [15:0] out_s1885;
wire  [15:0] out_s1886;
wire  [15:0] out_s1887;
wire  [15:0] out_s1888;
wire  [15:0] out_s1889;
wire  [15:0] out_s1890;
wire  [15:0] out_s1891;
wire  [15:0] out_s1892;
wire  [15:0] out_s1893;
wire  [15:0] out_s1894;
wire  [15:0] out_s1895;
wire  [15:0] out_s1896;
wire  [15:0] out_s1897;
wire  [15:0] out_s1898;
wire  [15:0] out_s1899;
wire  [15:0] out_s1900;
wire  [15:0] out_s1901;
wire  [15:0] out_s1902;
wire  [15:0] out_s1903;
wire  [15:0] out_s1904;
wire  [15:0] out_s1905;
wire  [15:0] out_s1906;
wire  [15:0] out_s1907;
wire  [15:0] out_s1908;
wire  [15:0] out_s1909;
wire  [15:0] out_s1910;
wire  [15:0] out_s1911;
wire  [15:0] out_s1912;
wire  [15:0] out_s1913;
wire  [15:0] out_s1914;
wire  [15:0] out_s1915;
wire  [15:0] out_s1916;
wire  [15:0] out_s1917;
wire  [15:0] out_s1918;
wire  [15:0] out_s1919;
wire  [15:0] out_s1920;
wire  [15:0] out_s1921;
wire  [15:0] out_s1922;
wire  [15:0] out_s1923;
wire  [15:0] out_s1924;
wire  [15:0] out_s1925;
wire  [15:0] out_s1926;
wire  [15:0] out_s1927;
wire  [15:0] out_s1928;
wire  [15:0] out_s1929;
wire  [15:0] out_s1930;
wire  [15:0] out_s1931;
wire  [15:0] out_s1932;
wire  [15:0] out_s1933;
wire  [15:0] out_s1934;
wire  [15:0] out_s1935;
wire  [15:0] out_s1936;
wire  [15:0] out_s1937;
wire  [15:0] out_s1938;
wire  [15:0] out_s1939;
wire  [15:0] out_s1940;
wire  [15:0] out_s1941;
wire  [15:0] out_s1942;
wire  [15:0] out_s1943;
wire  [15:0] out_s1944;
wire  [15:0] out_s1945;
wire  [15:0] out_s1946;
wire  [15:0] out_s1947;
wire  [15:0] out_s1948;
wire  [15:0] out_s1949;
wire  [15:0] out_s1950;
wire  [15:0] out_s1951;
wire  [15:0] out_s1952;
wire  [15:0] out_s1953;
wire  [15:0] out_s1954;
wire  [15:0] out_s1955;
wire  [15:0] out_s1956;
wire  [15:0] out_s1957;
wire  [15:0] out_s1958;
wire  [15:0] out_s1959;
wire  [15:0] out_s1960;
wire  [15:0] out_s1961;
wire  [15:0] out_s1962;
wire  [15:0] out_s1963;
wire  [15:0] out_s1964;
wire  [15:0] out_s1965;
wire  [15:0] out_s1966;
wire  [15:0] out_s1967;
wire  [15:0] out_s1968;
wire  [15:0] out_s1969;
wire  [15:0] out_s1970;
wire  [15:0] out_s1971;
wire  [15:0] out_s1972;
wire  [15:0] out_s1973;
wire  [15:0] out_s1974;
wire  [15:0] out_s1975;
wire  [15:0] out_s1976;
wire  [15:0] out_s1977;
wire  [15:0] out_s1978;
wire  [15:0] out_s1979;
wire  [15:0] out_s1980;
wire  [15:0] out_s1981;
wire  [15:0] out_s1982;
wire  [15:0] out_s1983;
wire  [15:0] out_s1984;
wire  [15:0] out_s1985;
wire  [15:0] out_s1986;
wire  [15:0] out_s1987;
wire  [15:0] out_s1988;
wire  [15:0] out_s1989;
wire  [15:0] out_s1990;
wire  [15:0] out_s1991;
wire  [15:0] out_s1992;
wire  [15:0] out_s1993;
wire  [15:0] out_s1994;
wire  [15:0] out_s1995;
wire  [15:0] out_s1996;
wire  [15:0] out_s1997;
wire  [15:0] out_s1998;
wire  [15:0] out_s1999;
wire  [15:0] out_s2000;
wire  [15:0] out_s2001;
wire  [15:0] out_s2002;
wire  [15:0] out_s2003;
wire  [15:0] out_s2004;
wire  [15:0] out_s2005;
wire  [15:0] out_s2006;
wire  [15:0] out_s2007;
wire  [15:0] out_s2008;
wire  [15:0] out_s2009;
wire  [15:0] out_s2010;
wire  [15:0] out_s2011;
wire  [15:0] out_s2012;
wire  [15:0] out_s2013;
wire  [15:0] out_s2014;
wire  [15:0] out_s2015;
wire  [15:0] out_s2016;
wire  [15:0] out_s2017;
wire  [15:0] out_s2018;
wire  [15:0] out_s2019;
wire  [15:0] out_s2020;
wire  [15:0] out_s2021;
wire  [15:0] out_s2022;
wire  [15:0] out_s2023;
wire  [15:0] out_s2024;
wire  [15:0] out_s2025;
wire  [15:0] out_s2026;
wire  [15:0] out_s2027;
wire  [15:0] out_s2028;
wire  [15:0] out_s2029;
wire  [15:0] out_s2030;
wire  [15:0] out_s2031;
wire  [15:0] out_s2032;
wire  [15:0] out_s2033;
wire  [15:0] out_s2034;
wire  [15:0] out_s2035;
wire  [15:0] out_s2036;
wire  [15:0] out_s2037;
wire  [15:0] out_s2038;
wire  [15:0] out_s2039;
wire  [15:0] out_s2040;
wire  [15:0] out_s2041;
wire  [15:0] out_s2042;
wire  [15:0] out_s2043;
wire  [15:0] out_s2044;
wire  [15:0] out_s2045;
wire  [15:0] out_s2046;
wire  [15:0] out_s2047;
wire  [15:0] out_s2048;
wire  [15:0] out_s2049;
wire  [15:0] out_s2050;
wire  [15:0] out_s2051;
wire  [15:0] out_s2052;
wire  [15:0] out_s2053;
wire  [15:0] out_s2054;
wire  [15:0] out_s2055;
wire  [15:0] out_s2056;
wire  [15:0] out_s2057;
wire  [15:0] out_s2058;
wire  [15:0] out_s2059;
wire  [15:0] out_s2060;
wire  [15:0] out_s2061;
wire  [15:0] out_s2062;
wire  [15:0] out_s2063;
wire  [15:0] out_s2064;
wire  [15:0] out_s2065;
wire  [15:0] out_s2066;
wire  [15:0] out_s2067;
wire  [15:0] out_s2068;
wire  [15:0] out_s2069;
wire  [15:0] out_s2070;
wire  [15:0] out_s2071;
wire  [15:0] out_s2072;
wire  [15:0] out_s2073;
wire  [15:0] out_s2074;
wire  [15:0] out_s2075;
wire  [15:0] out_s2076;
wire  [15:0] out_s2077;
wire  [15:0] out_s2078;
wire  [15:0] out_s2079;
wire  [15:0] out_s2080;
wire  [15:0] out_s2081;
wire  [15:0] out_s2082;
wire  [15:0] out_s2083;
wire  [15:0] out_s2084;
wire  [15:0] out_s2085;
wire  [15:0] out_s2086;
wire  [15:0] out_s2087;
wire  [15:0] out_s2088;
wire  [15:0] out_s2089;
wire  [15:0] out_s2090;
wire  [15:0] out_s2091;
wire  [15:0] out_s2092;
wire  [15:0] out_s2093;
wire  [15:0] out_s2094;
wire  [15:0] out_s2095;
wire  [15:0] out_s2096;
wire  [15:0] out_s2097;
wire  [15:0] out_s2098;
wire  [15:0] out_s2099;
wire  [15:0] out_s2100;
wire  [15:0] out_s2101;
wire  [15:0] out_s2102;
wire  [15:0] out_s2103;
wire  [15:0] out_s2104;
wire  [15:0] out_s2105;
wire  [15:0] out_s2106;
wire  [15:0] out_s2107;
wire  [15:0] out_s2108;
wire  [15:0] out_s2109;
wire  [15:0] out_s2110;
wire  [15:0] out_s2111;
wire  [15:0] out_s2112;
wire  [15:0] out_s2113;
wire  [15:0] out_s2114;
wire  [15:0] out_s2115;
wire  [15:0] out_s2116;
wire  [15:0] out_s2117;
wire  [15:0] out_s2118;
wire  [15:0] out_s2119;
wire  [15:0] out_s2120;
wire  [15:0] out_s2121;
wire  [15:0] out_s2122;
wire  [15:0] out_s2123;
wire  [15:0] out_s2124;
wire  [15:0] out_s2125;
wire  [15:0] out_s2126;
wire  [15:0] out_s2127;
wire  [15:0] out_s2128;
wire  [15:0] out_s2129;
wire  [15:0] out_s2130;
wire  [15:0] out_s2131;
wire  [15:0] out_s2132;
wire  [15:0] out_s2133;
wire  [15:0] out_s2134;
wire  [15:0] out_s2135;
wire  [15:0] out_s2136;
wire  [15:0] out_s2137;
wire  [15:0] out_s2138;
wire  [15:0] out_s2139;
wire  [15:0] out_s2140;
wire  [15:0] out_s2141;
wire  [15:0] out_s2142;
wire  [15:0] out_s2143;
wire  [15:0] out_s2144;
wire  [15:0] out_s2145;
wire  [15:0] out_s2146;
wire  [15:0] out_s2147;
wire  [15:0] out_s2148;
wire  [15:0] out_s2149;
wire  [15:0] out_s2150;
wire  [15:0] out_s2151;
wire  [15:0] out_s2152;
wire  [15:0] out_s2153;
wire  [15:0] out_s2154;
wire  [15:0] out_s2155;
wire  [15:0] out_s2156;
wire  [15:0] out_s2157;
wire  [15:0] out_s2158;
wire  [15:0] out_s2159;
wire  [15:0] out_s2160;
wire  [15:0] out_s2161;
wire  [15:0] out_s2162;
wire  [15:0] out_s2163;
wire  [15:0] out_s2164;
wire  [15:0] out_s2165;
wire  [15:0] out_s2166;
wire  [15:0] out_s2167;
wire  [15:0] out_s2168;
wire  [15:0] out_s2169;
wire  [15:0] out_s2170;
wire  [15:0] out_s2171;
wire  [15:0] out_s2172;
wire  [15:0] out_s2173;
wire  [15:0] out_s2174;
wire  [15:0] out_s2175;
wire  [15:0] out_s2176;
wire  [15:0] out_s2177;
wire  [15:0] out_s2178;
wire  [15:0] out_s2179;
wire  [15:0] out_s2180;
wire  [15:0] out_s2181;
wire  [15:0] out_s2182;
wire  [15:0] out_s2183;
wire  [15:0] out_s2184;
wire  [15:0] out_s2185;
wire  [15:0] out_s2186;
wire  [15:0] out_s2187;
wire  [15:0] out_s2188;
wire  [15:0] out_s2189;
wire  [15:0] out_s2190;
wire  [15:0] out_s2191;
wire  [15:0] out_s2192;
wire  [15:0] out_s2193;
wire  [15:0] out_s2194;
wire  [15:0] out_s2195;
wire  [15:0] out_s2196;
wire  [15:0] out_s2197;
wire  [15:0] out_s2198;
wire  [15:0] out_s2199;
wire  [15:0] out_s2200;
wire  [15:0] out_s2201;
wire  [15:0] out_s2202;
wire  [15:0] out_s2203;
wire  [15:0] out_s2204;
wire  [15:0] out_s2205;
wire  [15:0] out_s2206;
wire  [15:0] out_s2207;
wire  [15:0] out_s2208;
wire  [15:0] out_s2209;
wire  [15:0] out_s2210;
wire  [15:0] out_s2211;
wire  [15:0] out_s2212;
wire  [15:0] out_s2213;
wire  [15:0] out_s2214;
wire  [15:0] out_s2215;
wire  [15:0] out_s2216;
wire  [15:0] out_s2217;
wire  [15:0] out_s2218;
wire  [15:0] out_s2219;
wire  [15:0] out_s2220;
wire  [15:0] out_s2221;
wire  [15:0] out_s2222;
wire  [15:0] out_s2223;
wire  [15:0] out_s2224;
wire  [15:0] out_s2225;
wire  [15:0] out_s2226;
wire  [15:0] out_s2227;
wire  [15:0] out_s2228;
wire  [15:0] out_s2229;
wire  [15:0] out_s2230;
wire  [15:0] out_s2231;
wire  [15:0] out_s2232;
wire  [15:0] out_s2233;
wire  [15:0] out_s2234;
wire  [15:0] out_s2235;
wire  [15:0] out_s2236;
wire  [15:0] out_s2237;
wire  [15:0] out_s2238;
wire  [15:0] out_s2239;
wire  [15:0] out_s2240;
wire  [15:0] out_s2241;
wire  [15:0] out_s2242;
wire  [15:0] out_s2243;
wire  [15:0] out_s2244;
wire  [15:0] out_s2245;
wire  [15:0] out_s2246;
wire  [15:0] out_s2247;
wire  [15:0] out_s2248;
wire  [15:0] out_s2249;
wire  [15:0] out_s2250;
wire  [15:0] out_s2251;
wire  [15:0] out_s2252;
wire  [15:0] out_s2253;
wire  [15:0] out_s2254;
wire  [15:0] out_s2255;
wire  [15:0] out_s2256;
wire  [15:0] out_s2257;
wire  [15:0] out_s2258;
wire  [15:0] out_s2259;
wire  [15:0] out_s2260;
wire  [15:0] out_s2261;
wire  [15:0] out_s2262;
wire  [15:0] out_s2263;
wire  [15:0] out_s2264;
wire  [15:0] out_s2265;
wire  [15:0] out_s2266;
wire  [15:0] out_s2267;
wire  [15:0] out_s2268;
wire  [15:0] out_s2269;
wire  [15:0] out_s2270;
wire  [15:0] out_s2271;
wire  [15:0] out_s2272;
wire  [15:0] out_s2273;
wire  [15:0] out_s2274;
wire  [15:0] out_s2275;
wire  [15:0] out_s2276;
wire  [15:0] out_s2277;
wire  [15:0] out_s2278;
wire  [15:0] out_s2279;
wire  [15:0] out_s2280;
wire  [15:0] out_s2281;
wire  [15:0] out_s2282;
wire  [15:0] out_s2283;
wire  [15:0] out_s2284;
wire  [15:0] out_s2285;
wire  [15:0] out_s2286;
wire  [15:0] out_s2287;
wire  [15:0] out_s2288;
wire  [15:0] out_s2289;
wire  [15:0] out_s2290;
wire  [15:0] out_s2291;
wire  [15:0] out_s2292;
wire  [15:0] out_s2293;
wire  [15:0] out_s2294;
wire  [15:0] out_s2295;
wire  [15:0] out_s2296;
wire  [15:0] out_s2297;
wire  [15:0] out_s2298;
wire  [15:0] out_s2299;
wire  [15:0] out_s2300;
wire  [15:0] out_s2301;
wire  [15:0] out_s2302;
wire  [15:0] out_s2303;
wire  [15:0] out_s2304;
wire  [15:0] out_s2305;
wire  [15:0] out_s2306;
wire  [15:0] out_s2307;
wire  [15:0] out_s2308;
wire  [15:0] out_s2309;
wire  [15:0] out_s2310;
wire  [15:0] out_s2311;
wire  [15:0] out_s2312;
wire  [15:0] out_s2313;
wire  [15:0] out_s2314;
wire  [15:0] out_s2315;
wire  [15:0] out_s2316;
wire  [15:0] out_s2317;
wire  [15:0] out_s2318;
wire  [15:0] out_s2319;
wire  [15:0] out_s2320;
wire  [15:0] out_s2321;
wire  [15:0] out_s2322;
wire  [15:0] out_s2323;
wire  [15:0] out_s2324;
wire  [15:0] out_s2325;
wire  [15:0] out_s2326;
wire  [15:0] out_s2327;
wire  [15:0] out_s2328;
wire  [15:0] out_s2329;
wire  [15:0] out_s2330;
wire  [15:0] out_s2331;
wire  [15:0] out_s2332;
wire  [15:0] out_s2333;
wire  [15:0] out_s2334;
wire  [15:0] out_s2335;
wire  [15:0] out_s2336;
wire  [15:0] out_s2337;
wire  [15:0] out_s2338;
wire  [15:0] out_s2339;
wire  [15:0] out_s2340;
wire  [15:0] out_s2341;
wire  [15:0] out_s2342;
wire  [15:0] out_s2343;
wire  [15:0] out_s2344;
wire  [15:0] out_s2345;
wire  [15:0] out_s2346;
wire  [15:0] out_s2347;
wire  [15:0] out_s2348;
wire  [15:0] out_s2349;
wire  [15:0] out_s2350;
wire  [15:0] out_s2351;
wire  [15:0] out_s2352;
wire  [15:0] out_s2353;
wire  [15:0] out_s2354;
wire  [15:0] out_s2355;
wire  [15:0] out_s2356;
wire  [15:0] out_s2357;
wire  [15:0] out_s2358;
wire  [15:0] out_s2359;
wire  [15:0] out_s2360;
wire  [15:0] out_s2361;
wire  [15:0] out_s2362;
wire  [15:0] out_s2363;
wire  [15:0] out_s2364;
wire  [15:0] out_s2365;
wire  [15:0] out_s2366;
wire  [15:0] out_s2367;
wire  [15:0] out_s2368;
wire  [15:0] out_s2369;
wire  [15:0] out_s2370;
wire  [15:0] out_s2371;
wire  [15:0] out_s2372;
wire  [15:0] out_s2373;
wire  [15:0] out_s2374;
wire  [15:0] out_s2375;
wire  [15:0] out_s2376;
wire  [15:0] out_s2377;
wire  [15:0] out_s2378;
wire  [15:0] out_s2379;
wire  [15:0] out_s2380;
wire  [15:0] out_s2381;
wire  [15:0] out_s2382;
wire  [15:0] out_s2383;
wire  [15:0] out_s2384;
wire  [15:0] out_s2385;
wire  [15:0] out_s2386;
wire  [15:0] out_s2387;
wire  [15:0] out_s2388;
wire  [15:0] out_s2389;
wire  [15:0] out_s2390;
wire  [15:0] out_s2391;
wire  [15:0] out_s2392;
wire  [15:0] out_s2393;
wire  [15:0] out_s2394;
wire  [15:0] out_s2395;
wire  [15:0] out_s2396;
wire  [15:0] out_s2397;
wire  [15:0] out_s2398;
wire  [15:0] out_s2399;
wire  [15:0] out_s2400;
wire  [15:0] out_s2401;
wire  [15:0] out_s2402;
wire  [15:0] out_s2403;
wire  [15:0] out_s2404;
wire  [15:0] out_s2405;
wire  [15:0] out_s2406;
wire  [15:0] out_s2407;
wire  [15:0] out_s2408;
wire  [15:0] out_s2409;
wire  [15:0] out_s2410;
wire  [15:0] out_s2411;
wire  [15:0] out_s2412;
wire  [15:0] out_s2413;
wire  [15:0] out_s2414;
wire  [15:0] out_s2415;
wire  [15:0] out_s2416;
wire  [15:0] out_s2417;
wire  [15:0] out_s2418;
wire  [15:0] out_s2419;
wire  [15:0] out_s2420;
wire  [15:0] out_s2421;
wire  [15:0] out_s2422;
wire  [15:0] out_s2423;
wire  [15:0] out_s2424;
wire  [15:0] out_s2425;
wire  [15:0] out_s2426;
wire  [15:0] out_s2427;
wire  [15:0] out_s2428;
wire  [15:0] out_s2429;
wire  [15:0] out_s2430;
wire  [15:0] out_s2431;
wire  [15:0] out_s2432;
wire  [15:0] out_s2433;
wire  [15:0] out_s2434;
wire  [15:0] out_s2435;
wire  [15:0] out_s2436;
wire  [15:0] out_s2437;
wire  [15:0] out_s2438;
wire  [15:0] out_s2439;
wire  [15:0] out_s2440;
wire  [15:0] out_s2441;
wire  [15:0] out_s2442;
wire  [15:0] out_s2443;
wire  [15:0] out_s2444;
wire  [15:0] out_s2445;
wire  [15:0] out_s2446;
wire  [15:0] out_s2447;
wire  [15:0] out_s2448;
wire  [15:0] out_s2449;
wire  [15:0] out_s2450;
wire  [15:0] out_s2451;
wire  [15:0] out_s2452;
wire  [15:0] out_s2453;
wire  [15:0] out_s2454;
wire  [15:0] out_s2455;
wire  [15:0] out_s2456;
wire  [15:0] out_s2457;
wire  [15:0] out_s2458;
wire  [15:0] out_s2459;
wire  [15:0] out_s2460;
wire  [15:0] out_s2461;
wire  [15:0] out_s2462;
wire  [15:0] out_s2463;
wire  [15:0] out_s2464;
wire  [15:0] out_s2465;
wire  [15:0] out_s2466;
wire  [15:0] out_s2467;
wire  [15:0] out_s2468;
wire  [15:0] out_s2469;
wire  [15:0] out_s2470;
wire  [15:0] out_s2471;
wire  [15:0] out_s2472;
wire  [15:0] out_s2473;
wire  [15:0] out_s2474;
wire  [15:0] out_s2475;
wire  [15:0] out_s2476;
wire  [15:0] out_s2477;
wire  [15:0] out_s2478;
wire  [15:0] out_s2479;
wire  [15:0] out_s2480;
wire  [15:0] out_s2481;
wire  [15:0] out_s2482;
wire  [15:0] out_s2483;
wire  [15:0] out_s2484;
wire  [15:0] out_s2485;
wire  [15:0] out_s2486;
wire  [15:0] out_s2487;
wire  [15:0] out_s2488;
wire  [15:0] out_s2489;
wire  [15:0] out_s2490;
wire  [15:0] out_s2491;
wire  [15:0] out_s2492;
wire  [15:0] out_s2493;
wire  [15:0] out_s2494;
wire  [15:0] out_s2495;
wire  [15:0] out_s2496;
wire  [15:0] out_s2497;
wire  [15:0] out_s2498;
wire  [15:0] out_s2499;
wire  [15:0] out_s2500;
wire  [15:0] out_s2501;
wire  [15:0] out_s2502;
wire  [15:0] out_s2503;
wire  [15:0] out_s2504;
wire  [15:0] out_s2505;
wire  [15:0] out_s2506;
wire  [15:0] out_s2507;
wire  [15:0] out_s2508;
wire  [15:0] out_s2509;
wire  [15:0] out_s2510;
wire  [15:0] out_s2511;
wire  [15:0] out_s2512;
wire  [15:0] out_s2513;
wire  [15:0] out_s2514;
wire  [15:0] out_s2515;
wire  [15:0] out_s2516;
wire  [15:0] out_s2517;
wire  [15:0] out_s2518;
wire  [15:0] out_s2519;
wire  [15:0] out_s2520;
wire  [15:0] out_s2521;
wire  [15:0] out_s2522;
wire  [15:0] out_s2523;
wire  [15:0] out_s2524;
wire  [15:0] out_s2525;
wire  [15:0] out_s2526;
wire  [15:0] out_s2527;
wire  [15:0] out_s2528;
wire  [15:0] out_s2529;
wire  [15:0] out_s2530;
wire  [15:0] out_s2531;
wire  [15:0] out_s2532;
wire  [15:0] out_s2533;
wire  [15:0] out_s2534;
wire  [15:0] out_s2535;
wire  [15:0] out_s2536;
wire  [15:0] out_s2537;
wire  [15:0] out_s2538;
wire  [15:0] out_s2539;
wire  [15:0] out_s2540;
wire  [15:0] out_s2541;
wire  [15:0] out_s2542;
wire  [15:0] out_s2543;
wire  [15:0] out_s2544;
wire  [15:0] out_s2545;
wire  [15:0] out_s2546;
wire  [15:0] out_s2547;
wire  [15:0] out_s2548;
wire  [15:0] out_s2549;
wire  [15:0] out_s2550;
wire  [15:0] out_s2551;
wire  [15:0] out_s2552;
wire  [15:0] out_s2553;
wire  [15:0] out_s2554;
wire  [15:0] out_s2555;
wire  [15:0] out_s2556;
wire  [15:0] out_s2557;
wire  [15:0] out_s2558;
wire  [15:0] out_s2559;
wire  [15:0] out_s2560;
wire  [15:0] out_s2561;
wire  [15:0] out_s2562;
wire  [15:0] out_s2563;
wire  [15:0] out_s2564;
wire  [15:0] out_s2565;
wire  [15:0] out_s2566;
wire  [15:0] out_s2567;
wire  [15:0] out_s2568;
wire  [15:0] out_s2569;
wire  [15:0] out_s2570;
wire  [15:0] out_s2571;
wire  [15:0] out_s2572;
wire  [15:0] out_s2573;
wire  [15:0] out_s2574;
wire  [15:0] out_s2575;
wire  [15:0] out_s2576;
wire  [15:0] out_s2577;
wire  [15:0] out_s2578;
wire  [15:0] out_s2579;
wire  [15:0] out_s2580;
wire  [15:0] out_s2581;
wire  [15:0] out_s2582;
wire  [15:0] out_s2583;
wire  [15:0] out_s2584;
wire  [15:0] out_s2585;
wire  [15:0] out_s2586;
wire  [15:0] out_s2587;
wire  [15:0] out_s2588;
wire  [15:0] out_s2589;
wire  [15:0] out_s2590;
wire  [15:0] out_s2591;
wire  [15:0] out_s2592;
wire  [15:0] out_s2593;
wire  [15:0] out_s2594;
wire  [15:0] out_s2595;
wire  [15:0] out_s2596;
wire  [15:0] out_s2597;
wire  [15:0] out_s2598;
wire  [15:0] out_s2599;
wire  [15:0] out_s2600;
wire  [15:0] out_s2601;
wire  [15:0] out_s2602;
wire  [15:0] out_s2603;
wire  [15:0] out_s2604;
wire  [15:0] out_s2605;
wire  [15:0] out_s2606;
wire  [15:0] out_s2607;
wire  [15:0] out_s2608;
wire  [15:0] out_s2609;
wire  [15:0] out_s2610;
wire  [15:0] out_s2611;
wire  [15:0] out_s2612;
wire  [15:0] out_s2613;
wire  [15:0] out_s2614;
wire  [15:0] out_s2615;
wire  [15:0] out_s2616;
wire  [15:0] out_s2617;
wire  [15:0] out_s2618;
wire  [15:0] out_s2619;
wire  [15:0] out_s2620;
wire  [15:0] out_s2621;
wire  [15:0] out_s2622;
wire  [15:0] out_s2623;
wire  [15:0] out_s2624;
wire  [15:0] out_s2625;
wire  [15:0] out_s2626;
wire  [15:0] out_s2627;
wire  [15:0] out_s2628;
wire  [15:0] out_s2629;
wire  [15:0] out_s2630;
wire  [15:0] out_s2631;
wire  [15:0] out_s2632;
wire  [15:0] out_s2633;
wire  [15:0] out_s2634;
wire  [15:0] out_s2635;
wire  [15:0] out_s2636;
wire  [15:0] out_s2637;
wire  [15:0] out_s2638;
wire  [15:0] out_s2639;
wire  [15:0] out_s2640;
wire  [15:0] out_s2641;
wire  [15:0] out_s2642;
wire  [15:0] out_s2643;
wire  [15:0] out_s2644;
wire  [15:0] out_s2645;
wire  [15:0] out_s2646;
wire  [15:0] out_s2647;
wire  [15:0] out_s2648;
wire  [15:0] out_s2649;
wire  [15:0] out_s2650;
wire  [15:0] out_s2651;
wire  [15:0] out_s2652;
wire  [15:0] out_s2653;
wire  [15:0] out_s2654;
wire  [15:0] out_s2655;
wire  [15:0] out_s2656;
wire  [15:0] out_s2657;
wire  [15:0] out_s2658;
wire  [15:0] out_s2659;
wire  [15:0] out_s2660;
wire  [15:0] out_s2661;
wire  [15:0] out_s2662;
wire  [15:0] out_s2663;
wire  [15:0] out_s2664;
wire  [15:0] out_s2665;
wire  [15:0] out_s2666;
wire  [15:0] out_s2667;
wire  [15:0] out_s2668;
wire  [15:0] out_s2669;
wire  [15:0] out_s2670;
wire  [15:0] out_s2671;
wire  [15:0] out_s2672;
wire  [15:0] out_s2673;
wire  [15:0] out_s2674;
wire  [15:0] out_s2675;
wire  [15:0] out_s2676;
wire  [15:0] out_s2677;
wire  [15:0] out_s2678;
wire  [15:0] out_s2679;
wire  [15:0] out_s2680;
wire  [15:0] out_s2681;
wire  [15:0] out_s2682;
wire  [15:0] out_s2683;
wire  [15:0] out_s2684;
wire  [15:0] out_s2685;
wire  [15:0] out_s2686;
wire  [15:0] out_s2687;
wire  [15:0] out_s2688;
wire  [15:0] out_s2689;
wire  [15:0] out_s2690;
wire  [15:0] out_s2691;
wire  [15:0] out_s2692;
wire  [15:0] out_s2693;
wire  [15:0] out_s2694;
wire  [15:0] out_s2695;
wire  [15:0] out_s2696;
wire  [15:0] out_s2697;
wire  [15:0] out_s2698;
wire  [15:0] out_s2699;
wire  [15:0] out_s2700;
wire  [15:0] out_s2701;
wire  [15:0] out_s2702;
wire  [15:0] out_s2703;
wire  [15:0] out_s2704;
wire  [15:0] out_s2705;
wire  [15:0] out_s2706;
wire  [15:0] out_s2707;
wire  [15:0] out_s2708;
wire  [15:0] out_s2709;
wire  [15:0] out_s2710;
wire  [15:0] out_s2711;
wire  [15:0] out_s2712;
wire  [15:0] out_s2713;
wire  [15:0] out_s2714;
wire  [15:0] out_s2715;
wire  [15:0] out_s2716;
wire  [15:0] out_s2717;
wire  [15:0] out_s2718;
wire  [15:0] out_s2719;
wire  [15:0] out_s2720;
wire  [15:0] out_s2721;
wire  [15:0] out_s2722;
wire  [15:0] out_s2723;
wire  [15:0] out_s2724;
wire  [15:0] out_s2725;
wire  [15:0] out_s2726;
wire  [15:0] out_s2727;
wire  [15:0] out_s2728;
wire  [15:0] out_s2729;
wire  [15:0] out_s2730;
wire  [15:0] out_s2731;
wire  [15:0] out_s2732;
wire  [15:0] out_s2733;
wire  [15:0] out_s2734;
wire  [15:0] out_s2735;
wire  [15:0] out_s2736;
wire  [15:0] out_s2737;
wire  [15:0] out_s2738;
wire  [15:0] out_s2739;
wire  [15:0] out_s2740;
wire  [15:0] out_s2741;
wire  [15:0] out_s2742;
wire  [15:0] out_s2743;
wire  [15:0] out_s2744;
wire  [15:0] out_s2745;
wire  [15:0] out_s2746;
wire  [15:0] out_s2747;
wire  [15:0] out_s2748;
wire  [15:0] out_s2749;
wire  [15:0] out_s2750;
wire  [15:0] out_s2751;
wire  [15:0] out_s2752;
wire  [15:0] out_s2753;
wire  [15:0] out_s2754;
wire  [15:0] out_s2755;
wire  [15:0] out_s2756;
wire  [15:0] out_s2757;
wire  [15:0] out_s2758;
wire  [15:0] out_s2759;
wire  [15:0] out_s2760;
wire  [15:0] out_s2761;
wire  [15:0] out_s2762;
wire  [15:0] out_s2763;
wire  [15:0] out_s2764;
wire  [15:0] out_s2765;
wire  [15:0] out_s2766;
wire  [15:0] out_s2767;
wire  [15:0] out_s2768;
wire  [15:0] out_s2769;
wire  [15:0] out_s2770;
wire  [15:0] out_s2771;
wire  [15:0] out_s2772;
wire  [15:0] out_s2773;
wire  [15:0] out_s2774;
wire  [15:0] out_s2775;
wire  [15:0] out_s2776;
wire  [15:0] out_s2777;
wire  [15:0] out_s2778;
wire  [15:0] out_s2779;
wire  [15:0] out_s2780;
wire  [15:0] out_s2781;
wire  [15:0] out_s2782;
wire  [15:0] out_s2783;
wire  [15:0] out_s2784;
wire  [15:0] out_s2785;
wire  [15:0] out_s2786;
wire  [15:0] out_s2787;
wire  [15:0] out_s2788;
wire  [15:0] out_s2789;
wire  [15:0] out_s2790;
wire  [15:0] out_s2791;
wire  [15:0] out_s2792;
wire  [15:0] out_s2793;
wire  [15:0] out_s2794;
wire  [15:0] out_s2795;
wire  [15:0] out_s2796;
wire  [15:0] out_s2797;
wire  [15:0] out_s2798;
wire  [15:0] out_s2799;
wire  [15:0] out_s2800;
wire  [15:0] out_s2801;
wire  [15:0] out_s2802;
wire  [15:0] out_s2803;
wire  [15:0] out_s2804;
wire  [15:0] out_s2805;
wire  [15:0] out_s2806;
wire  [15:0] out_s2807;
wire  [15:0] out_s2808;
wire  [15:0] out_s2809;
wire  [15:0] out_s2810;
wire  [15:0] out_s2811;
wire  [15:0] out_s2812;
wire  [15:0] out_s2813;
wire  [15:0] out_s2814;
wire  [15:0] out_s2815;
wire  [15:0] out_s2816;
wire  [15:0] out_s2817;
wire  [15:0] out_s2818;
wire  [15:0] out_s2819;
wire  [15:0] out_s2820;
wire  [15:0] out_s2821;
wire  [15:0] out_s2822;
wire  [15:0] out_s2823;
wire  [15:0] out_s2824;
wire  [15:0] out_s2825;
wire  [15:0] out_s2826;
wire  [15:0] out_s2827;
wire  [15:0] out_s2828;
wire  [15:0] out_s2829;
wire  [15:0] out_s2830;
wire  [15:0] out_s2831;
wire  [15:0] out_s2832;
wire  [15:0] out_s2833;
wire  [15:0] out_s2834;
wire  [15:0] out_s2835;
wire  [15:0] out_s2836;
wire  [15:0] out_s2837;
wire  [15:0] out_s2838;
wire  [15:0] out_s2839;
wire  [15:0] out_s2840;
wire  [15:0] out_s2841;
wire  [15:0] out_s2842;
wire  [15:0] out_s2843;
wire  [15:0] out_s2844;
wire  [15:0] out_s2845;
wire  [15:0] out_s2846;
wire  [15:0] out_s2847;
wire  [15:0] out_s2848;
wire  [15:0] out_s2849;
wire  [15:0] out_s2850;
wire  [15:0] out_s2851;
wire  [15:0] out_s2852;
wire  [15:0] out_s2853;
wire  [15:0] out_s2854;
wire  [15:0] out_s2855;
wire  [15:0] out_s2856;
wire  [15:0] out_s2857;
wire  [15:0] out_s2858;
wire  [15:0] out_s2859;
wire  [15:0] out_s2860;
wire  [15:0] out_s2861;
wire  [15:0] out_s2862;
wire  [15:0] out_s2863;
wire  [15:0] out_s2864;
wire  [15:0] out_s2865;
wire  [15:0] out_s2866;
wire  [15:0] out_s2867;
wire  [15:0] out_s2868;
wire  [15:0] out_s2869;
wire  [15:0] out_s2870;
wire  [15:0] out_s2871;
wire  [15:0] out_s2872;
wire  [15:0] out_s2873;
wire  [15:0] out_s2874;
wire  [15:0] out_s2875;
wire  [15:0] out_s2876;
wire  [15:0] out_s2877;
wire  [15:0] out_s2878;
wire  [15:0] out_s2879;
wire  [15:0] out_s2880;
wire  [15:0] out_s2881;
wire  [15:0] out_s2882;
wire  [15:0] out_s2883;
wire  [15:0] out_s2884;
wire  [15:0] out_s2885;
wire  [15:0] out_s2886;
wire  [15:0] out_s2887;
wire  [15:0] out_s2888;
wire  [15:0] out_s2889;
wire  [15:0] out_s2890;
wire  [15:0] out_s2891;
wire  [15:0] out_s2892;
wire  [15:0] out_s2893;
wire  [15:0] out_s2894;
wire  [15:0] out_s2895;
wire  [15:0] out_s2896;
wire  [15:0] out_s2897;
wire  [15:0] out_s2898;
wire  [15:0] out_s2899;
wire  [15:0] out_s2900;
wire  [15:0] out_s2901;
wire  [15:0] out_s2902;
wire  [15:0] out_s2903;
wire  [15:0] out_s2904;
wire  [15:0] out_s2905;
wire  [15:0] out_s2906;
wire  [15:0] out_s2907;
wire  [15:0] out_s2908;
wire  [15:0] out_s2909;
wire  [15:0] out_s2910;
wire  [15:0] out_s2911;
wire  [15:0] out_s2912;
wire  [15:0] out_s2913;
wire  [15:0] out_s2914;
wire  [15:0] out_s2915;
wire  [15:0] out_s2916;
wire  [15:0] out_s2917;
wire  [15:0] out_s2918;
wire  [15:0] out_s2919;
wire  [15:0] out_s2920;
wire  [15:0] out_s2921;
wire  [15:0] out_s2922;
wire  [15:0] out_s2923;
wire  [15:0] out_s2924;
wire  [15:0] out_s2925;
wire  [15:0] out_s2926;
wire  [15:0] out_s2927;
wire  [15:0] out_s2928;
wire  [15:0] out_s2929;
wire  [15:0] out_s2930;
wire  [15:0] out_s2931;
wire  [15:0] out_s2932;
wire  [15:0] out_s2933;
wire  [15:0] out_s2934;
wire  [15:0] out_s2935;
wire  [15:0] out_s2936;
wire  [15:0] out_s2937;
wire  [15:0] out_s2938;
wire  [15:0] out_s2939;
wire  [15:0] out_s2940;
wire  [15:0] out_s2941;
wire  [15:0] out_s2942;
wire  [15:0] out_s2943;
wire  [15:0] out_s2944;
wire  [15:0] out_s2945;
wire  [15:0] out_s2946;
wire  [15:0] out_s2947;
wire  [15:0] out_s2948;
wire  [15:0] out_s2949;
wire  [15:0] out_s2950;
wire  [15:0] out_s2951;
wire  [15:0] out_s2952;
wire  [15:0] out_s2953;
wire  [15:0] out_s2954;
wire  [15:0] out_s2955;
wire  [15:0] out_s2956;
wire  [15:0] out_s2957;
wire  [15:0] out_s2958;
wire  [15:0] out_s2959;
wire  [15:0] out_s2960;
wire  [15:0] out_s2961;
wire  [15:0] out_s2962;
wire  [15:0] out_s2963;
wire  [15:0] out_s2964;
wire  [15:0] out_s2965;
wire  [15:0] out_s2966;
wire  [15:0] out_s2967;
wire  [15:0] out_s2968;
wire  [15:0] out_s2969;
wire  [15:0] out_s2970;
wire  [15:0] out_s2971;
wire  [15:0] out_s2972;
wire  [15:0] out_s2973;
wire  [15:0] out_s2974;
wire  [15:0] out_s2975;
wire  [15:0] out_s2976;
wire  [15:0] out_s2977;
wire  [15:0] out_s2978;
wire  [15:0] out_s2979;
wire  [15:0] out_s2980;
wire  [15:0] out_s2981;
wire  [15:0] out_s2982;
wire  [15:0] out_s2983;
wire  [15:0] out_s2984;
wire  [15:0] out_s2985;
wire  [15:0] out_s2986;
wire  [15:0] out_s2987;
wire  [15:0] out_s2988;
wire  [15:0] out_s2989;
wire  [15:0] out_s2990;
wire  [15:0] out_s2991;
wire  [15:0] out_s2992;
wire  [15:0] out_s2993;
wire  [15:0] out_s2994;
wire  [15:0] out_s2995;
wire  [15:0] out_s2996;
wire  [15:0] out_s2997;
wire  [15:0] out_s2998;
wire  [15:0] out_s2999;
wire  [15:0] out_s3000;
wire  [15:0] out_s3001;
wire  [15:0] out_s3002;
wire  [15:0] out_s3003;
wire  [15:0] out_s3004;
wire  [15:0] out_s3005;
wire  [15:0] out_s3006;
wire  [15:0] out_s3007;
wire  [15:0] out_s3008;
wire  [15:0] out_s3009;
wire  [15:0] out_s3010;
wire  [15:0] out_s3011;
wire  [15:0] out_s3012;
wire  [15:0] out_s3013;
wire  [15:0] out_s3014;
wire  [15:0] out_s3015;
wire  [15:0] out_s3016;
wire  [15:0] out_s3017;
wire  [15:0] out_s3018;
wire  [15:0] out_s3019;
wire  [15:0] out_s3020;
wire  [15:0] out_s3021;
wire  [15:0] out_s3022;
wire  [15:0] out_s3023;
wire  [15:0] out_s3024;
wire  [15:0] out_s3025;
wire  [15:0] out_s3026;
wire  [15:0] out_s3027;
wire  [15:0] out_s3028;
wire  [15:0] out_s3029;
wire  [15:0] out_s3030;
wire  [15:0] out_s3031;
wire  [15:0] out_s3032;
wire  [15:0] out_s3033;
wire  [15:0] out_s3034;
wire  [15:0] out_s3035;
wire  [15:0] out_s3036;
wire  [15:0] out_s3037;
wire  [15:0] out_s3038;
wire  [15:0] out_s3039;
wire  [15:0] out_s3040;
wire  [15:0] out_s3041;
wire  [15:0] out_s3042;
wire  [15:0] out_s3043;
wire  [15:0] out_s3044;
wire  [15:0] out_s3045;
wire  [15:0] out_s3046;
wire  [15:0] out_s3047;
wire  [15:0] out_s3048;
wire  [15:0] out_s3049;
wire  [15:0] out_s3050;
wire  [15:0] out_s3051;
wire  [15:0] out_s3052;
wire  [15:0] out_s3053;
wire  [15:0] out_s3054;
wire  [15:0] out_s3055;
wire  [15:0] out_s3056;
wire  [15:0] out_s3057;
wire  [15:0] out_s3058;
wire  [15:0] out_s3059;
wire  [15:0] out_s3060;
wire  [15:0] out_s3061;
wire  [15:0] out_s3062;
wire  [15:0] out_s3063;
wire  [15:0] out_s3064;
wire  [15:0] out_s3065;
wire  [15:0] out_s3066;
wire  [15:0] out_s3067;
wire  [15:0] out_s3068;
wire  [15:0] out_s3069;
wire  [15:0] out_s3070;
wire  [15:0] out_s3071;
wire  [15:0] out_s3072;
wire  [15:0] out_s3073;
wire  [15:0] out_s3074;
wire  [15:0] out_s3075;
wire  [15:0] out_s3076;
wire  [15:0] out_s3077;
wire  [15:0] out_s3078;
wire  [15:0] out_s3079;
wire  [15:0] out_s3080;
wire  [15:0] out_s3081;
wire  [15:0] out_s3082;
wire  [15:0] out_s3083;
wire  [15:0] out_s3084;
wire  [15:0] out_s3085;
wire  [15:0] out_s3086;
wire  [15:0] out_s3087;
wire  [15:0] out_s3088;
wire  [15:0] out_s3089;
wire  [15:0] out_s3090;
wire  [15:0] out_s3091;
wire  [15:0] out_s3092;
wire  [15:0] out_s3093;
wire  [15:0] out_s3094;
wire  [15:0] out_s3095;
wire  [15:0] out_s3096;
wire  [15:0] out_s3097;
wire  [15:0] out_s3098;
wire  [15:0] out_s3099;
wire  [15:0] out_s3100;
wire  [15:0] out_s3101;
wire  [15:0] out_s3102;
wire  [15:0] out_s3103;
wire  [15:0] out_s3104;
wire  [15:0] out_s3105;
wire  [15:0] out_s3106;
wire  [15:0] out_s3107;
wire  [15:0] out_s3108;
wire  [15:0] out_s3109;
wire  [15:0] out_s3110;
wire  [15:0] out_s3111;
wire  [15:0] out_s3112;
wire  [15:0] out_s3113;
wire  [15:0] out_s3114;
wire  [15:0] out_s3115;
wire  [15:0] out_s3116;
wire  [15:0] out_s3117;
wire  [15:0] out_s3118;
wire  [15:0] out_s3119;
wire  [15:0] out_s3120;
wire  [15:0] out_s3121;
wire  [15:0] out_s3122;
wire  [15:0] out_s3123;
wire  [15:0] out_s3124;
wire  [15:0] out_s3125;
wire  [15:0] out_s3126;
wire  [15:0] out_s3127;
wire  [15:0] out_s3128;
wire  [15:0] out_s3129;
wire  [15:0] out_s3130;
wire  [15:0] out_s3131;
wire  [15:0] out_s3132;
wire  [15:0] out_s3133;
wire  [15:0] out_s3134;
wire  [15:0] out_s3135;
wire  [15:0] out_s3136;
wire  [15:0] out_s3137;
wire  [15:0] out_s3138;
wire  [15:0] out_s3139;
wire  [15:0] out_s3140;
wire  [15:0] out_s3141;
wire  [15:0] out_s3142;
wire  [15:0] out_s3143;
wire  [15:0] out_s3144;
wire  [15:0] out_s3145;
wire  [15:0] out_s3146;
wire  [15:0] out_s3147;
wire  [15:0] out_s3148;
wire  [15:0] out_s3149;
wire  [15:0] out_s3150;
wire  [15:0] out_s3151;
wire  [15:0] out_s3152;
wire  [15:0] out_s3153;
wire  [15:0] out_s3154;
wire  [15:0] out_s3155;
wire  [15:0] out_s3156;
wire  [15:0] out_s3157;
wire  [15:0] out_s3158;
wire  [15:0] out_s3159;
wire  [15:0] out_s3160;
wire  [15:0] out_s3161;
wire  [15:0] out_s3162;
wire  [15:0] out_s3163;
wire  [15:0] out_s3164;
wire  [15:0] out_s3165;
wire  [15:0] out_s3166;
wire  [15:0] out_s3167;
wire  [15:0] out_s3168;
wire  [15:0] out_s3169;
wire  [15:0] out_s3170;
wire  [15:0] out_s3171;
wire  [15:0] out_s3172;
wire  [15:0] out_s3173;
wire  [15:0] out_s3174;
wire  [15:0] out_s3175;
wire  [15:0] out_s3176;
wire  [15:0] out_s3177;
wire  [15:0] out_s3178;
wire  [15:0] out_s3179;
wire  [15:0] out_s3180;
wire  [15:0] out_s3181;
wire  [15:0] out_s3182;
wire  [15:0] out_s3183;
wire  [15:0] out_s3184;
wire  [15:0] out_s3185;
wire  [15:0] out_s3186;
wire  [15:0] out_s3187;
wire  [15:0] out_s3188;
wire  [15:0] out_s3189;
wire  [15:0] out_s3190;
wire  [15:0] out_s3191;
wire  [15:0] out_s3192;
wire  [15:0] out_s3193;
wire  [15:0] out_s3194;
wire  [15:0] out_s3195;
wire  [15:0] out_s3196;
wire  [15:0] out_s3197;
wire  [15:0] out_s3198;
wire  [15:0] out_s3199;
wire  [15:0] out_s3200;
wire  [15:0] out_s3201;
wire  [15:0] out_s3202;
wire  [15:0] out_s3203;
wire  [15:0] out_s3204;
wire  [15:0] out_s3205;
wire  [15:0] out_s3206;
wire  [15:0] out_s3207;
wire  [15:0] out_s3208;
wire  [15:0] out_s3209;
wire  [15:0] out_s3210;
wire  [15:0] out_s3211;
wire  [15:0] out_s3212;
wire  [15:0] out_s3213;
wire  [15:0] out_s3214;
wire  [15:0] out_s3215;
wire  [15:0] out_s3216;
wire  [15:0] out_s3217;
wire  [15:0] out_s3218;
wire  [15:0] out_s3219;
wire  [15:0] out_s3220;
wire  [15:0] out_s3221;
wire  [15:0] out_s3222;
wire  [15:0] out_s3223;
wire  [15:0] out_s3224;
wire  [15:0] out_s3225;
wire  [15:0] out_s3226;
wire  [15:0] out_s3227;
wire  [15:0] out_s3228;
wire  [15:0] out_s3229;
wire  [15:0] out_s3230;
wire  [15:0] out_s3231;
wire  [15:0] out_s3232;
wire  [15:0] out_s3233;
wire  [15:0] out_s3234;
wire  [15:0] out_s3235;
wire  [15:0] out_s3236;
wire  [15:0] out_s3237;
wire  [15:0] out_s3238;
wire  [15:0] out_s3239;
wire  [15:0] out_s3240;
wire  [15:0] out_s3241;
wire  [15:0] out_s3242;
wire  [15:0] out_s3243;
wire  [15:0] out_s3244;
wire  [15:0] out_s3245;
wire  [15:0] out_s3246;
wire  [15:0] out_s3247;
wire  [15:0] out_s3248;
wire  [15:0] out_s3249;
wire  [15:0] out_s3250;
wire  [15:0] out_s3251;
wire  [15:0] out_s3252;
wire  [15:0] out_s3253;
wire  [15:0] out_s3254;
wire  [15:0] out_s3255;
wire  [15:0] out_s3256;
wire  [15:0] out_s3257;
wire  [15:0] out_s3258;
wire  [15:0] out_s3259;
wire  [15:0] out_s3260;
wire  [15:0] out_s3261;
wire  [15:0] out_s3262;
wire  [15:0] out_s3263;
wire  [15:0] out_s3264;
wire  [15:0] out_s3265;
wire  [15:0] out_s3266;
wire  [15:0] out_s3267;
wire  [15:0] out_s3268;
wire  [15:0] out_s3269;
wire  [15:0] out_s3270;
wire  [15:0] out_s3271;
wire  [15:0] out_s3272;
wire  [15:0] out_s3273;
wire  [15:0] out_s3274;
wire  [15:0] out_s3275;
wire  [15:0] out_s3276;
wire  [15:0] out_s3277;
wire  [15:0] out_s3278;
wire  [15:0] out_s3279;
wire  [15:0] out_s3280;
wire  [15:0] out_s3281;
wire  [15:0] out_s3282;
wire  [15:0] out_s3283;
wire  [15:0] out_s3284;
wire  [15:0] out_s3285;
wire  [15:0] out_s3286;
wire  [15:0] out_s3287;
wire  [15:0] out_s3288;
wire  [15:0] out_s3289;
wire  [15:0] out_s3290;
wire  [15:0] out_s3291;
wire  [15:0] out_s3292;
wire  [15:0] out_s3293;
wire  [15:0] out_s3294;
wire  [15:0] out_s3295;
wire  [15:0] out_s3296;
wire  [15:0] out_s3297;
wire  [15:0] out_s3298;
wire  [15:0] out_s3299;
wire  [15:0] out_s3300;
wire  [15:0] out_s3301;
wire  [15:0] out_s3302;
wire  [15:0] out_s3303;
wire  [15:0] out_s3304;
wire  [15:0] out_s3305;
wire  [15:0] out_s3306;
wire  [15:0] out_s3307;
wire  [15:0] out_s3308;
wire  [15:0] out_s3309;
wire  [15:0] out_s3310;
wire  [15:0] out_s3311;
wire  [15:0] out_s3312;
wire  [15:0] out_s3313;
wire  [15:0] out_s3314;
wire  [15:0] out_s3315;
wire  [15:0] out_s3316;
wire  [15:0] out_s3317;
wire  [15:0] out_s3318;
wire  [15:0] out_s3319;
wire  [15:0] out_s3320;
wire  [15:0] out_s3321;
wire  [15:0] out_s3322;
wire  [15:0] out_s3323;
wire  [15:0] out_s3324;
wire  [15:0] out_s3325;
wire  [15:0] out_s3326;
wire  [15:0] out_s3327;
wire  [15:0] out_s3328;
wire  [15:0] out_s3329;
wire  [15:0] out_s3330;
wire  [15:0] out_s3331;
wire  [15:0] out_s3332;
wire  [15:0] out_s3333;
wire  [15:0] out_s3334;
wire  [15:0] out_s3335;
wire  [15:0] out_s3336;
wire  [15:0] out_s3337;
wire  [15:0] out_s3338;
wire  [15:0] out_s3339;
wire  [15:0] out_s3340;
wire  [15:0] out_s3341;
wire  [15:0] out_s3342;
wire  [15:0] out_s3343;
wire  [15:0] out_s3344;
wire  [15:0] out_s3345;
wire  [15:0] out_s3346;
wire  [15:0] out_s3347;
wire  [15:0] out_s3348;
wire  [15:0] out_s3349;
wire  [15:0] out_s3350;
wire  [15:0] out_s3351;
wire  [15:0] out_s3352;
wire  [15:0] out_s3353;
wire  [15:0] out_s3354;
wire  [15:0] out_s3355;
wire  [15:0] out_s3356;
wire  [15:0] out_s3357;
wire  [15:0] out_s3358;
wire  [15:0] out_s3359;
wire  [15:0] out_s3360;
wire  [15:0] out_s3361;
wire  [15:0] out_s3362;
wire  [15:0] out_s3363;
wire  [15:0] out_s3364;
wire  [15:0] out_s3365;
wire  [15:0] out_s3366;
wire  [15:0] out_s3367;
wire  [15:0] out_s3368;
wire  [15:0] out_s3369;
wire  [15:0] out_s3370;
wire  [15:0] out_s3371;
wire  [15:0] out_s3372;
wire  [15:0] out_s3373;
wire  [15:0] out_s3374;
wire  [15:0] out_s3375;
wire  [15:0] out_s3376;
wire  [15:0] out_s3377;
wire  [15:0] out_s3378;
wire  [15:0] out_s3379;
wire  [15:0] out_s3380;
wire  [15:0] out_s3381;
wire  [15:0] out_s3382;
wire  [15:0] out_s3383;
wire  [15:0] out_s3384;
wire  [15:0] out_s3385;
wire  [15:0] out_s3386;
wire  [15:0] out_s3387;
wire  [15:0] out_s3388;
wire  [15:0] out_s3389;
wire  [15:0] out_s3390;
wire  [15:0] out_s3391;
wire  [15:0] out_s3392;
wire  [15:0] out_s3393;
wire  [15:0] out_s3394;
wire  [15:0] out_s3395;
wire  [15:0] out_s3396;
wire  [15:0] out_s3397;
wire  [15:0] out_s3398;
wire  [15:0] out_s3399;
wire  [15:0] out_s3400;
wire  [15:0] out_s3401;
wire  [15:0] out_s3402;
wire  [15:0] out_s3403;
wire  [15:0] out_s3404;
wire  [15:0] out_s3405;
wire  [15:0] out_s3406;
wire  [15:0] out_s3407;
wire  [15:0] out_s3408;
wire  [15:0] out_s3409;
wire  [15:0] out_s3410;
wire  [15:0] out_s3411;
wire  [15:0] out_s3412;
wire  [15:0] out_s3413;
wire  [15:0] out_s3414;
wire  [15:0] out_s3415;
wire  [15:0] out_s3416;
wire  [15:0] out_s3417;
wire  [15:0] out_s3418;
wire  [15:0] out_s3419;
wire  [15:0] out_s3420;
wire  [15:0] out_s3421;
wire  [15:0] out_s3422;
wire  [15:0] out_s3423;
wire  [15:0] out_s3424;
wire  [15:0] out_s3425;
wire  [15:0] out_s3426;
wire  [15:0] out_s3427;
wire  [15:0] out_s3428;
wire  [15:0] out_s3429;
wire  [15:0] out_s3430;
wire  [15:0] out_s3431;
wire  [15:0] out_s3432;
wire  [15:0] out_s3433;
wire  [15:0] out_s3434;
wire  [15:0] out_s3435;
wire  [15:0] out_s3436;
wire  [15:0] out_s3437;
wire  [15:0] out_s3438;
wire  [15:0] out_s3439;
wire  [15:0] out_s3440;
wire  [15:0] out_s3441;
wire  [15:0] out_s3442;
wire  [15:0] out_s3443;
wire  [15:0] out_s3444;
wire  [15:0] out_s3445;
wire  [15:0] out_s3446;
wire  [15:0] out_s3447;
wire  [15:0] out_s3448;
wire  [15:0] out_s3449;
wire  [15:0] out_s3450;
wire  [15:0] out_s3451;
wire  [15:0] out_s3452;
wire  [15:0] out_s3453;
wire  [15:0] out_s3454;
wire  [15:0] out_s3455;
wire  [15:0] out_s3456;
wire  [15:0] out_s3457;
wire  [15:0] out_s3458;
wire  [15:0] out_s3459;
wire  [15:0] out_s3460;
wire  [15:0] out_s3461;
wire  [15:0] out_s3462;
wire  [15:0] out_s3463;
wire  [15:0] out_s3464;
wire  [15:0] out_s3465;
wire  [15:0] out_s3466;
wire  [15:0] out_s3467;
wire  [15:0] out_s3468;
wire  [15:0] out_s3469;
wire  [15:0] out_s3470;
wire  [15:0] out_s3471;
wire  [15:0] out_s3472;
wire  [15:0] out_s3473;
wire  [15:0] out_s3474;
wire  [15:0] out_s3475;
wire  [15:0] out_s3476;
wire  [15:0] out_s3477;
wire  [15:0] out_s3478;
wire  [15:0] out_s3479;
wire  [15:0] out_s3480;
wire  [15:0] out_s3481;
wire  [15:0] out_s3482;
wire  [15:0] out_s3483;
wire  [15:0] out_s3484;
wire  [15:0] out_s3485;
wire  [15:0] out_s3486;
wire  [15:0] out_s3487;
wire  [15:0] out_s3488;
wire  [15:0] out_s3489;
wire  [15:0] out_s3490;
wire  [15:0] out_s3491;
wire  [15:0] out_s3492;
wire  [15:0] out_s3493;
wire  [15:0] out_s3494;
wire  [15:0] out_s3495;
wire  [15:0] out_s3496;
wire  [15:0] out_s3497;
wire  [15:0] out_s3498;
wire  [15:0] out_s3499;
wire  [15:0] out_s3500;
wire  [15:0] out_s3501;
wire  [15:0] out_s3502;
wire  [15:0] out_s3503;
wire  [15:0] out_s3504;
wire  [15:0] out_s3505;
wire  [15:0] out_s3506;
wire  [15:0] out_s3507;
wire  [15:0] out_s3508;
wire  [15:0] out_s3509;
wire  [15:0] out_s3510;
wire  [15:0] out_s3511;
wire  [15:0] out_s3512;
wire  [15:0] out_s3513;
wire  [15:0] out_s3514;
wire  [15:0] out_s3515;
wire  [15:0] out_s3516;
wire  [15:0] out_s3517;
wire  [15:0] out_s3518;
wire  [15:0] out_s3519;
wire  [15:0] out_s3520;
wire  [15:0] out_s3521;
wire  [15:0] out_s3522;
wire  [15:0] out_s3523;
wire  [15:0] out_s3524;
wire  [15:0] out_s3525;
wire  [15:0] out_s3526;
wire  [15:0] out_s3527;
wire  [15:0] out_s3528;
wire  [15:0] out_s3529;
wire  [15:0] out_s3530;
wire  [15:0] out_s3531;
wire  [15:0] out_s3532;
wire  [15:0] out_s3533;
wire  [15:0] out_s3534;
wire  [15:0] out_s3535;
wire  [15:0] out_s3536;
wire  [15:0] out_s3537;
wire  [15:0] out_s3538;
wire  [15:0] out_s3539;
wire  [15:0] out_s3540;
wire  [15:0] out_s3541;
wire  [15:0] out_s3542;
wire  [15:0] out_s3543;
wire  [15:0] out_s3544;
wire  [15:0] out_s3545;
wire  [15:0] out_s3546;
wire  [15:0] out_s3547;
wire  [15:0] out_s3548;
wire  [15:0] out_s3549;
wire  [15:0] out_s3550;
wire  [15:0] out_s3551;
wire  [15:0] out_s3552;
wire  [15:0] out_s3553;
wire  [15:0] out_s3554;
wire  [15:0] out_s3555;
wire  [15:0] out_s3556;
wire  [15:0] out_s3557;
wire  [15:0] out_s3558;
wire  [15:0] out_s3559;
wire  [15:0] out_s3560;
wire  [15:0] out_s3561;
wire  [15:0] out_s3562;
wire  [15:0] out_s3563;
wire  [15:0] out_s3564;
wire  [15:0] out_s3565;
wire  [15:0] out_s3566;
wire  [15:0] out_s3567;
wire  [15:0] out_s3568;
wire  [15:0] out_s3569;
wire  [15:0] out_s3570;
wire  [15:0] out_s3571;
wire  [15:0] out_s3572;
wire  [15:0] out_s3573;
wire  [15:0] out_s3574;
wire  [15:0] out_s3575;
wire  [15:0] out_s3576;
wire  [15:0] out_s3577;
wire  [15:0] out_s3578;
wire  [15:0] out_s3579;
wire  [15:0] out_s3580;
wire  [15:0] out_s3581;
wire  [15:0] out_s3582;
wire  [15:0] out_s3583;
wire  [15:0] out_s3584;
wire  [15:0] out_s3585;
wire  [15:0] out_s3586;
wire  [15:0] out_s3587;
wire  [15:0] out_s3588;
wire  [15:0] out_s3589;
wire  [15:0] out_s3590;
wire  [15:0] out_s3591;
wire  [15:0] out_s3592;
wire  [15:0] out_s3593;
wire  [15:0] out_s3594;
wire  [15:0] out_s3595;
wire  [15:0] out_s3596;
wire  [15:0] out_s3597;
wire  [15:0] out_s3598;
wire  [15:0] out_s3599;
wire  [15:0] out_s3600;
wire  [15:0] out_s3601;
wire  [15:0] out_s3602;
wire  [15:0] out_s3603;
wire  [15:0] out_s3604;
wire  [15:0] out_s3605;
wire  [15:0] out_s3606;
wire  [15:0] out_s3607;
wire  [15:0] out_s3608;
wire  [15:0] out_s3609;
wire  [15:0] out_s3610;
wire  [15:0] out_s3611;
wire  [15:0] out_s3612;
wire  [15:0] out_s3613;
wire  [15:0] out_s3614;
wire  [15:0] out_s3615;
wire  [15:0] out_s3616;
wire  [15:0] out_s3617;
wire  [15:0] out_s3618;
wire  [15:0] out_s3619;
wire  [15:0] out_s3620;
wire  [15:0] out_s3621;
wire  [15:0] out_s3622;
wire  [15:0] out_s3623;
wire  [15:0] out_s3624;
wire  [15:0] out_s3625;
wire  [15:0] out_s3626;
wire  [15:0] out_s3627;
wire  [15:0] out_s3628;
wire  [15:0] out_s3629;
wire  [15:0] out_s3630;
wire  [15:0] out_s3631;
wire  [15:0] out_s3632;
wire  [15:0] out_s3633;
wire  [15:0] out_s3634;
wire  [15:0] out_s3635;
wire  [15:0] out_s3636;
wire  [15:0] out_s3637;
wire  [15:0] out_s3638;
wire  [15:0] out_s3639;
wire  [15:0] out_s3640;
wire  [15:0] out_s3641;
wire  [15:0] out_s3642;
wire  [15:0] out_s3643;
wire  [15:0] out_s3644;
wire  [15:0] out_s3645;
wire  [15:0] out_s3646;
wire  [15:0] out_s3647;
wire  [15:0] out_s3648;
wire  [15:0] out_s3649;
wire  [15:0] out_s3650;
wire  [15:0] out_s3651;
wire  [15:0] out_s3652;
wire  [15:0] out_s3653;
wire  [15:0] out_s3654;
wire  [15:0] out_s3655;
wire  [15:0] out_s3656;
wire  [15:0] out_s3657;
wire  [15:0] out_s3658;
wire  [15:0] out_s3659;
wire  [15:0] out_s3660;
wire  [15:0] out_s3661;
wire  [15:0] out_s3662;
wire  [15:0] out_s3663;
wire  [15:0] out_s3664;
wire  [15:0] out_s3665;
wire  [15:0] out_s3666;
wire  [15:0] out_s3667;
wire  [15:0] out_s3668;
wire  [15:0] out_s3669;
wire  [15:0] out_s3670;
wire  [15:0] out_s3671;
wire  [15:0] out_s3672;
wire  [15:0] out_s3673;
wire  [15:0] out_s3674;
wire  [15:0] out_s3675;
wire  [15:0] out_s3676;
wire  [15:0] out_s3677;
wire  [15:0] out_s3678;
wire  [15:0] out_s3679;
wire  [15:0] out_s3680;
wire  [15:0] out_s3681;
wire  [15:0] out_s3682;
wire  [15:0] out_s3683;
wire  [15:0] out_s3684;
wire  [15:0] out_s3685;
wire  [15:0] out_s3686;
wire  [15:0] out_s3687;
wire  [15:0] out_s3688;
wire  [15:0] out_s3689;
wire  [15:0] out_s3690;
wire  [15:0] out_s3691;
wire  [15:0] out_s3692;
wire  [15:0] out_s3693;
wire  [15:0] out_s3694;
wire  [15:0] out_s3695;
wire  [15:0] out_s3696;
wire  [15:0] out_s3697;
wire  [15:0] out_s3698;
wire  [15:0] out_s3699;
wire  [15:0] out_s3700;
wire  [15:0] out_s3701;
wire  [15:0] out_s3702;
wire  [15:0] out_s3703;
wire  [15:0] out_s3704;
wire  [15:0] out_s3705;
wire  [15:0] out_s3706;
wire  [15:0] out_s3707;
wire  [15:0] out_s3708;
wire  [15:0] out_s3709;
wire  [15:0] out_s3710;
wire  [15:0] out_s3711;
wire  [15:0] out_s3712;
wire  [15:0] out_s3713;
wire  [15:0] out_s3714;
wire  [15:0] out_s3715;
wire  [15:0] out_s3716;
wire  [15:0] out_s3717;
wire  [15:0] out_s3718;
wire  [15:0] out_s3719;
wire  [15:0] out_s3720;
wire  [15:0] out_s3721;
wire  [15:0] out_s3722;
wire  [15:0] out_s3723;
wire  [15:0] out_s3724;
wire  [15:0] out_s3725;
wire  [15:0] out_s3726;
wire  [15:0] out_s3727;
wire  [15:0] out_s3728;
wire  [15:0] out_s3729;
wire  [15:0] out_s3730;
wire  [15:0] out_s3731;
wire  [15:0] out_s3732;
wire  [15:0] out_s3733;
wire  [15:0] out_s3734;
wire  [15:0] out_s3735;
wire  [15:0] out_s3736;
wire  [15:0] out_s3737;
wire  [15:0] out_s3738;
wire  [15:0] out_s3739;
wire  [15:0] out_s3740;
wire  [15:0] out_s3741;
wire  [15:0] out_s3742;
wire  [15:0] out_s3743;
wire  [15:0] out_s3744;
wire  [15:0] out_s3745;
wire  [15:0] out_s3746;
wire  [15:0] out_s3747;
wire  [15:0] out_s3748;
wire  [15:0] out_s3749;
wire  [15:0] out_s3750;
wire  [15:0] out_s3751;
wire  [15:0] out_s3752;
wire  [15:0] out_s3753;
wire  [15:0] out_s3754;
wire  [15:0] out_s3755;
wire  [15:0] out_s3756;
wire  [15:0] out_s3757;
wire  [15:0] out_s3758;
wire  [15:0] out_s3759;
wire  [15:0] out_s3760;
wire  [15:0] out_s3761;
wire  [15:0] out_s3762;
wire  [15:0] out_s3763;
wire  [15:0] out_s3764;
wire  [15:0] out_s3765;
wire  [15:0] out_s3766;
wire  [15:0] out_s3767;
wire  [15:0] out_s3768;
wire  [15:0] out_s3769;
wire  [15:0] out_s3770;
wire  [15:0] out_s3771;
wire  [15:0] out_s3772;
wire  [15:0] out_s3773;
wire  [15:0] out_s3774;
wire  [15:0] out_s3775;
wire  [15:0] out_s3776;
wire  [15:0] out_s3777;
wire  [15:0] out_s3778;
wire  [15:0] out_s3779;
wire  [15:0] out_s3780;
wire  [15:0] out_s3781;
wire  [15:0] out_s3782;
wire  [15:0] out_s3783;
wire  [15:0] out_s3784;
wire  [15:0] out_s3785;
wire  [15:0] out_s3786;
wire  [15:0] out_s3787;
wire  [15:0] out_s3788;
wire  [15:0] out_s3789;
wire  [15:0] out_s3790;
wire  [15:0] out_s3791;
wire  [15:0] out_s3792;
wire  [15:0] out_s3793;
wire  [15:0] out_s3794;
wire  [15:0] out_s3795;
wire  [15:0] out_s3796;
wire  [15:0] out_s3797;
wire  [15:0] out_s3798;
wire  [15:0] out_s3799;
wire  [15:0] out_s3800;
wire  [15:0] out_s3801;
wire  [15:0] out_s3802;
wire  [15:0] out_s3803;
wire  [15:0] out_s3804;
wire  [15:0] out_s3805;
wire  [15:0] out_s3806;
wire  [15:0] out_s3807;
wire  [15:0] out_s3808;
wire  [15:0] out_s3809;
wire  [15:0] out_s3810;
wire  [15:0] out_s3811;
wire  [15:0] out_s3812;
wire  [15:0] out_s3813;
wire  [15:0] out_s3814;
wire  [15:0] out_s3815;
wire  [15:0] out_s3816;
wire  [15:0] out_s3817;
wire  [15:0] out_s3818;
wire  [15:0] out_s3819;
wire  [15:0] out_s3820;
wire  [15:0] out_s3821;
wire  [15:0] out_s3822;
wire  [15:0] out_s3823;
wire  [15:0] out_s3824;
wire  [15:0] out_s3825;
wire  [15:0] out_s3826;
wire  [15:0] out_s3827;
wire  [15:0] out_s3828;
wire  [15:0] out_s3829;
wire  [15:0] out_s3830;
wire  [15:0] out_s3831;
wire  [15:0] out_s3832;
wire  [15:0] out_s3833;
wire  [15:0] out_s3834;
wire  [15:0] out_s3835;
wire  [15:0] out_s3836;
wire  [15:0] out_s3837;
wire  [15:0] out_s3838;
wire  [15:0] out_s3839;
wire  [15:0] out_s3840;
wire  [15:0] out_s3841;
wire  [15:0] out_s3842;
wire  [15:0] out_s3843;
wire  [15:0] out_s3844;
wire  [15:0] out_s3845;
wire  [15:0] out_s3846;
wire  [15:0] out_s3847;
wire  [15:0] out_s3848;
wire  [15:0] out_s3849;
wire  [15:0] out_s3850;
wire  [15:0] out_s3851;
wire  [15:0] out_s3852;
wire  [15:0] out_s3853;
wire  [15:0] out_s3854;
wire  [15:0] out_s3855;
wire  [15:0] out_s3856;
wire  [15:0] out_s3857;
wire  [15:0] out_s3858;
wire  [15:0] out_s3859;
wire  [15:0] out_s3860;
wire  [15:0] out_s3861;
wire  [15:0] out_s3862;
wire  [15:0] out_s3863;
wire  [15:0] out_s3864;
wire  [15:0] out_s3865;
wire  [15:0] out_s3866;
wire  [15:0] out_s3867;
wire  [15:0] out_s3868;
wire  [15:0] out_s3869;
wire  [15:0] out_s3870;
wire  [15:0] out_s3871;
wire  [15:0] out_s3872;
wire  [15:0] out_s3873;
wire  [15:0] out_s3874;
wire  [15:0] out_s3875;
wire  [15:0] out_s3876;
wire  [15:0] out_s3877;
wire  [15:0] out_s3878;
wire  [15:0] out_s3879;
wire  [15:0] out_s3880;
wire  [15:0] out_s3881;
wire  [15:0] out_s3882;
wire  [15:0] out_s3883;
wire  [15:0] out_s3884;
wire  [15:0] out_s3885;
wire  [15:0] out_s3886;
wire  [15:0] out_s3887;
wire  [15:0] out_s3888;
wire  [15:0] out_s3889;
wire  [15:0] out_s3890;
wire  [15:0] out_s3891;
wire  [15:0] out_s3892;
wire  [15:0] out_s3893;
wire  [15:0] out_s3894;
wire  [15:0] out_s3895;
wire  [15:0] out_s3896;
wire  [15:0] out_s3897;
wire  [15:0] out_s3898;
wire  [15:0] out_s3899;
wire  [15:0] out_s3900;
wire  [15:0] out_s3901;
wire  [15:0] out_s3902;
wire  [15:0] out_s3903;
wire  [15:0] out_s3904;
wire  [15:0] out_s3905;
wire  [15:0] out_s3906;
wire  [15:0] out_s3907;
wire  [15:0] out_s3908;
wire  [15:0] out_s3909;
wire  [15:0] out_s3910;
wire  [15:0] out_s3911;
wire  [15:0] out_s3912;
wire  [15:0] out_s3913;
wire  [15:0] out_s3914;
wire  [15:0] out_s3915;
wire  [15:0] out_s3916;
wire  [15:0] out_s3917;
wire  [15:0] out_s3918;
wire  [15:0] out_s3919;
wire  [15:0] out_s3920;
wire  [15:0] out_s3921;
wire  [15:0] out_s3922;
wire  [15:0] out_s3923;
wire  [15:0] out_s3924;
wire  [15:0] out_s3925;
wire  [15:0] out_s3926;
wire  [15:0] out_s3927;
wire  [15:0] out_s3928;
wire  [15:0] out_s3929;
wire  [15:0] out_s3930;
wire  [15:0] out_s3931;
wire  [15:0] out_s3932;
wire  [15:0] out_s3933;
wire  [15:0] out_s3934;
wire  [15:0] out_s3935;
wire  [15:0] out_s3936;
wire  [15:0] out_s3937;
wire  [15:0] out_s3938;
wire  [15:0] out_s3939;
wire  [15:0] out_s3940;
wire  [15:0] out_s3941;
wire  [15:0] out_s3942;
wire  [15:0] out_s3943;
wire  [15:0] out_s3944;
wire  [15:0] out_s3945;
wire  [15:0] out_s3946;
wire  [15:0] out_s3947;
wire  [15:0] out_s3948;
wire  [15:0] out_s3949;
wire  [15:0] out_s3950;
wire  [15:0] out_s3951;
wire  [15:0] out_s3952;
wire  [15:0] out_s3953;
wire  [15:0] out_s3954;
wire  [15:0] out_s3955;
wire  [15:0] out_s3956;
wire  [15:0] out_s3957;
wire  [15:0] out_s3958;
wire  [15:0] out_s3959;
wire  [15:0] out_s3960;
wire  [15:0] out_s3961;
wire  [15:0] out_s3962;
wire  [15:0] out_s3963;
wire  [15:0] out_s3964;
wire  [15:0] out_s3965;
wire  [15:0] out_s3966;
wire  [15:0] out_s3967;
wire  [15:0] out_s3968;
wire  [15:0] out_s3969;
wire  [15:0] out_s3970;
wire  [15:0] out_s3971;
wire  [15:0] out_s3972;
wire  [15:0] out_s3973;
wire  [15:0] out_s3974;
wire  [15:0] out_s3975;
wire  [15:0] out_s3976;
wire  [15:0] out_s3977;
wire  [15:0] out_s3978;
wire  [15:0] out_s3979;
wire  [15:0] out_s3980;
wire  [15:0] out_s3981;
wire  [15:0] out_s3982;
wire  [15:0] out_s3983;
wire  [15:0] out_s3984;
wire  [15:0] out_s3985;
wire  [15:0] out_s3986;
wire  [15:0] out_s3987;
wire  [15:0] out_s3988;
wire  [15:0] out_s3989;
wire  [15:0] out_s3990;
wire  [15:0] out_s3991;
wire  [15:0] out_s3992;
wire  [15:0] out_s3993;
wire  [15:0] out_s3994;
wire  [15:0] out_s3995;
wire  [15:0] out_s3996;
wire  [15:0] out_s3997;
wire  [15:0] out_s3998;
wire  [15:0] out_s3999;
wire  [15:0] out_s4000;
wire  [15:0] out_s4001;
wire  [15:0] out_s4002;
wire  [15:0] out_s4003;
wire  [15:0] out_s4004;
wire  [15:0] out_s4005;
wire  [15:0] out_s4006;
wire  [15:0] out_s4007;
wire  [15:0] out_s4008;
wire  [15:0] out_s4009;
wire  [15:0] out_s4010;
wire  [15:0] out_s4011;
wire  [15:0] out_s4012;
wire  [15:0] out_s4013;
wire  [15:0] out_s4014;
wire  [15:0] out_s4015;
wire  [15:0] out_s4016;
wire  [15:0] out_s4017;
wire  [15:0] out_s4018;
wire  [15:0] out_s4019;
wire  [15:0] out_s4020;
wire  [15:0] out_s4021;
wire  [15:0] out_s4022;
wire  [15:0] out_s4023;
wire  [15:0] out_s4024;
wire  [15:0] out_s4025;
wire  [15:0] out_s4026;
wire  [15:0] out_s4027;
wire  [15:0] out_s4028;
wire  [15:0] out_s4029;
wire  [15:0] out_s4030;
wire  [15:0] out_s4031;
wire  [15:0] out_s4032;
wire  [15:0] out_s4033;
wire  [15:0] out_s4034;
wire  [15:0] out_s4035;
wire  [15:0] out_s4036;
wire  [15:0] out_s4037;
wire  [15:0] out_s4038;
wire  [15:0] out_s4039;
wire  [15:0] out_s4040;
wire  [15:0] out_s4041;
wire  [15:0] out_s4042;
wire  [15:0] out_s4043;
wire  [15:0] out_s4044;
wire  [15:0] out_s4045;
wire  [15:0] out_s4046;
wire  [15:0] out_s4047;
wire  [15:0] out_s4048;
wire  [15:0] out_s4049;
wire  [15:0] out_s4050;
wire  [15:0] out_s4051;
wire  [15:0] out_s4052;
wire  [15:0] out_s4053;
wire  [15:0] out_s4054;
wire  [15:0] out_s4055;
wire  [15:0] out_s4056;
wire  [15:0] out_s4057;
wire  [15:0] out_s4058;
wire  [15:0] out_s4059;
wire  [15:0] out_s4060;
wire  [15:0] out_s4061;
wire  [15:0] out_s4062;
wire  [15:0] out_s4063;
wire  [15:0] out_s4064;
wire  [15:0] out_s4065;
wire  [15:0] out_s4066;
wire  [15:0] out_s4067;
wire  [15:0] out_s4068;
wire  [15:0] out_s4069;
wire  [15:0] out_s4070;
wire  [15:0] out_s4071;
wire  [15:0] out_s4072;
wire  [15:0] out_s4073;
wire  [15:0] out_s4074;
wire  [15:0] out_s4075;
wire  [15:0] out_s4076;
wire  [15:0] out_s4077;
wire  [15:0] out_s4078;
wire  [15:0] out_s4079;
wire  [15:0] out_s4080;
wire  [15:0] out_s4081;
wire  [15:0] out_s4082;
wire  [15:0] out_s4083;
wire  [15:0] out_s4084;
wire  [15:0] out_s4085;
wire  [15:0] out_s4086;
wire  [15:0] out_s4087;
wire  [15:0] out_s4088;
wire  [15:0] out_s4089;
wire  [15:0] out_s4090;
wire  [15:0] out_s4091;
wire  [15:0] out_s4092;
wire  [15:0] out_s4093;
wire  [15:0] out_s4094;
wire  [15:0] out_s4095;

wire  [15:0] out_e0;
wire  [15:0] out_e1;
wire  [15:0] out_e2;
wire  [15:0] out_e3;
wire  [15:0] out_e4;
wire  [15:0] out_e5;
wire  [15:0] out_e6;
wire  [15:0] out_e7;
wire  [15:0] out_e8;
wire  [15:0] out_e9;
wire  [15:0] out_e10;
wire  [15:0] out_e11;
wire  [15:0] out_e12;
wire  [15:0] out_e13;
wire  [15:0] out_e14;
wire  [15:0] out_e15;
wire  [15:0] out_e16;
wire  [15:0] out_e17;
wire  [15:0] out_e18;
wire  [15:0] out_e19;
wire  [15:0] out_e20;
wire  [15:0] out_e21;
wire  [15:0] out_e22;
wire  [15:0] out_e23;
wire  [15:0] out_e24;
wire  [15:0] out_e25;
wire  [15:0] out_e26;
wire  [15:0] out_e27;
wire  [15:0] out_e28;
wire  [15:0] out_e29;
wire  [15:0] out_e30;
wire  [15:0] out_e31;
wire  [15:0] out_e32;
wire  [15:0] out_e33;
wire  [15:0] out_e34;
wire  [15:0] out_e35;
wire  [15:0] out_e36;
wire  [15:0] out_e37;
wire  [15:0] out_e38;
wire  [15:0] out_e39;
wire  [15:0] out_e40;
wire  [15:0] out_e41;
wire  [15:0] out_e42;
wire  [15:0] out_e43;
wire  [15:0] out_e44;
wire  [15:0] out_e45;
wire  [15:0] out_e46;
wire  [15:0] out_e47;
wire  [15:0] out_e48;
wire  [15:0] out_e49;
wire  [15:0] out_e50;
wire  [15:0] out_e51;
wire  [15:0] out_e52;
wire  [15:0] out_e53;
wire  [15:0] out_e54;
wire  [15:0] out_e55;
wire  [15:0] out_e56;
wire  [15:0] out_e57;
wire  [15:0] out_e58;
wire  [15:0] out_e59;
wire  [15:0] out_e60;
wire  [15:0] out_e61;
wire  [15:0] out_e62;
wire  [15:0] out_e63;
wire  [15:0] out_e64;
wire  [15:0] out_e65;
wire  [15:0] out_e66;
wire  [15:0] out_e67;
wire  [15:0] out_e68;
wire  [15:0] out_e69;
wire  [15:0] out_e70;
wire  [15:0] out_e71;
wire  [15:0] out_e72;
wire  [15:0] out_e73;
wire  [15:0] out_e74;
wire  [15:0] out_e75;
wire  [15:0] out_e76;
wire  [15:0] out_e77;
wire  [15:0] out_e78;
wire  [15:0] out_e79;
wire  [15:0] out_e80;
wire  [15:0] out_e81;
wire  [15:0] out_e82;
wire  [15:0] out_e83;
wire  [15:0] out_e84;
wire  [15:0] out_e85;
wire  [15:0] out_e86;
wire  [15:0] out_e87;
wire  [15:0] out_e88;
wire  [15:0] out_e89;
wire  [15:0] out_e90;
wire  [15:0] out_e91;
wire  [15:0] out_e92;
wire  [15:0] out_e93;
wire  [15:0] out_e94;
wire  [15:0] out_e95;
wire  [15:0] out_e96;
wire  [15:0] out_e97;
wire  [15:0] out_e98;
wire  [15:0] out_e99;
wire  [15:0] out_e100;
wire  [15:0] out_e101;
wire  [15:0] out_e102;
wire  [15:0] out_e103;
wire  [15:0] out_e104;
wire  [15:0] out_e105;
wire  [15:0] out_e106;
wire  [15:0] out_e107;
wire  [15:0] out_e108;
wire  [15:0] out_e109;
wire  [15:0] out_e110;
wire  [15:0] out_e111;
wire  [15:0] out_e112;
wire  [15:0] out_e113;
wire  [15:0] out_e114;
wire  [15:0] out_e115;
wire  [15:0] out_e116;
wire  [15:0] out_e117;
wire  [15:0] out_e118;
wire  [15:0] out_e119;
wire  [15:0] out_e120;
wire  [15:0] out_e121;
wire  [15:0] out_e122;
wire  [15:0] out_e123;
wire  [15:0] out_e124;
wire  [15:0] out_e125;
wire  [15:0] out_e126;
wire  [15:0] out_e127;
wire  [15:0] out_e128;
wire  [15:0] out_e129;
wire  [15:0] out_e130;
wire  [15:0] out_e131;
wire  [15:0] out_e132;
wire  [15:0] out_e133;
wire  [15:0] out_e134;
wire  [15:0] out_e135;
wire  [15:0] out_e136;
wire  [15:0] out_e137;
wire  [15:0] out_e138;
wire  [15:0] out_e139;
wire  [15:0] out_e140;
wire  [15:0] out_e141;
wire  [15:0] out_e142;
wire  [15:0] out_e143;
wire  [15:0] out_e144;
wire  [15:0] out_e145;
wire  [15:0] out_e146;
wire  [15:0] out_e147;
wire  [15:0] out_e148;
wire  [15:0] out_e149;
wire  [15:0] out_e150;
wire  [15:0] out_e151;
wire  [15:0] out_e152;
wire  [15:0] out_e153;
wire  [15:0] out_e154;
wire  [15:0] out_e155;
wire  [15:0] out_e156;
wire  [15:0] out_e157;
wire  [15:0] out_e158;
wire  [15:0] out_e159;
wire  [15:0] out_e160;
wire  [15:0] out_e161;
wire  [15:0] out_e162;
wire  [15:0] out_e163;
wire  [15:0] out_e164;
wire  [15:0] out_e165;
wire  [15:0] out_e166;
wire  [15:0] out_e167;
wire  [15:0] out_e168;
wire  [15:0] out_e169;
wire  [15:0] out_e170;
wire  [15:0] out_e171;
wire  [15:0] out_e172;
wire  [15:0] out_e173;
wire  [15:0] out_e174;
wire  [15:0] out_e175;
wire  [15:0] out_e176;
wire  [15:0] out_e177;
wire  [15:0] out_e178;
wire  [15:0] out_e179;
wire  [15:0] out_e180;
wire  [15:0] out_e181;
wire  [15:0] out_e182;
wire  [15:0] out_e183;
wire  [15:0] out_e184;
wire  [15:0] out_e185;
wire  [15:0] out_e186;
wire  [15:0] out_e187;
wire  [15:0] out_e188;
wire  [15:0] out_e189;
wire  [15:0] out_e190;
wire  [15:0] out_e191;
wire  [15:0] out_e192;
wire  [15:0] out_e193;
wire  [15:0] out_e194;
wire  [15:0] out_e195;
wire  [15:0] out_e196;
wire  [15:0] out_e197;
wire  [15:0] out_e198;
wire  [15:0] out_e199;
wire  [15:0] out_e200;
wire  [15:0] out_e201;
wire  [15:0] out_e202;
wire  [15:0] out_e203;
wire  [15:0] out_e204;
wire  [15:0] out_e205;
wire  [15:0] out_e206;
wire  [15:0] out_e207;
wire  [15:0] out_e208;
wire  [15:0] out_e209;
wire  [15:0] out_e210;
wire  [15:0] out_e211;
wire  [15:0] out_e212;
wire  [15:0] out_e213;
wire  [15:0] out_e214;
wire  [15:0] out_e215;
wire  [15:0] out_e216;
wire  [15:0] out_e217;
wire  [15:0] out_e218;
wire  [15:0] out_e219;
wire  [15:0] out_e220;
wire  [15:0] out_e221;
wire  [15:0] out_e222;
wire  [15:0] out_e223;
wire  [15:0] out_e224;
wire  [15:0] out_e225;
wire  [15:0] out_e226;
wire  [15:0] out_e227;
wire  [15:0] out_e228;
wire  [15:0] out_e229;
wire  [15:0] out_e230;
wire  [15:0] out_e231;
wire  [15:0] out_e232;
wire  [15:0] out_e233;
wire  [15:0] out_e234;
wire  [15:0] out_e235;
wire  [15:0] out_e236;
wire  [15:0] out_e237;
wire  [15:0] out_e238;
wire  [15:0] out_e239;
wire  [15:0] out_e240;
wire  [15:0] out_e241;
wire  [15:0] out_e242;
wire  [15:0] out_e243;
wire  [15:0] out_e244;
wire  [15:0] out_e245;
wire  [15:0] out_e246;
wire  [15:0] out_e247;
wire  [15:0] out_e248;
wire  [15:0] out_e249;
wire  [15:0] out_e250;
wire  [15:0] out_e251;
wire  [15:0] out_e252;
wire  [15:0] out_e253;
wire  [15:0] out_e254;
wire  [15:0] out_e255;
wire  [15:0] out_e256;
wire  [15:0] out_e257;
wire  [15:0] out_e258;
wire  [15:0] out_e259;
wire  [15:0] out_e260;
wire  [15:0] out_e261;
wire  [15:0] out_e262;
wire  [15:0] out_e263;
wire  [15:0] out_e264;
wire  [15:0] out_e265;
wire  [15:0] out_e266;
wire  [15:0] out_e267;
wire  [15:0] out_e268;
wire  [15:0] out_e269;
wire  [15:0] out_e270;
wire  [15:0] out_e271;
wire  [15:0] out_e272;
wire  [15:0] out_e273;
wire  [15:0] out_e274;
wire  [15:0] out_e275;
wire  [15:0] out_e276;
wire  [15:0] out_e277;
wire  [15:0] out_e278;
wire  [15:0] out_e279;
wire  [15:0] out_e280;
wire  [15:0] out_e281;
wire  [15:0] out_e282;
wire  [15:0] out_e283;
wire  [15:0] out_e284;
wire  [15:0] out_e285;
wire  [15:0] out_e286;
wire  [15:0] out_e287;
wire  [15:0] out_e288;
wire  [15:0] out_e289;
wire  [15:0] out_e290;
wire  [15:0] out_e291;
wire  [15:0] out_e292;
wire  [15:0] out_e293;
wire  [15:0] out_e294;
wire  [15:0] out_e295;
wire  [15:0] out_e296;
wire  [15:0] out_e297;
wire  [15:0] out_e298;
wire  [15:0] out_e299;
wire  [15:0] out_e300;
wire  [15:0] out_e301;
wire  [15:0] out_e302;
wire  [15:0] out_e303;
wire  [15:0] out_e304;
wire  [15:0] out_e305;
wire  [15:0] out_e306;
wire  [15:0] out_e307;
wire  [15:0] out_e308;
wire  [15:0] out_e309;
wire  [15:0] out_e310;
wire  [15:0] out_e311;
wire  [15:0] out_e312;
wire  [15:0] out_e313;
wire  [15:0] out_e314;
wire  [15:0] out_e315;
wire  [15:0] out_e316;
wire  [15:0] out_e317;
wire  [15:0] out_e318;
wire  [15:0] out_e319;
wire  [15:0] out_e320;
wire  [15:0] out_e321;
wire  [15:0] out_e322;
wire  [15:0] out_e323;
wire  [15:0] out_e324;
wire  [15:0] out_e325;
wire  [15:0] out_e326;
wire  [15:0] out_e327;
wire  [15:0] out_e328;
wire  [15:0] out_e329;
wire  [15:0] out_e330;
wire  [15:0] out_e331;
wire  [15:0] out_e332;
wire  [15:0] out_e333;
wire  [15:0] out_e334;
wire  [15:0] out_e335;
wire  [15:0] out_e336;
wire  [15:0] out_e337;
wire  [15:0] out_e338;
wire  [15:0] out_e339;
wire  [15:0] out_e340;
wire  [15:0] out_e341;
wire  [15:0] out_e342;
wire  [15:0] out_e343;
wire  [15:0] out_e344;
wire  [15:0] out_e345;
wire  [15:0] out_e346;
wire  [15:0] out_e347;
wire  [15:0] out_e348;
wire  [15:0] out_e349;
wire  [15:0] out_e350;
wire  [15:0] out_e351;
wire  [15:0] out_e352;
wire  [15:0] out_e353;
wire  [15:0] out_e354;
wire  [15:0] out_e355;
wire  [15:0] out_e356;
wire  [15:0] out_e357;
wire  [15:0] out_e358;
wire  [15:0] out_e359;
wire  [15:0] out_e360;
wire  [15:0] out_e361;
wire  [15:0] out_e362;
wire  [15:0] out_e363;
wire  [15:0] out_e364;
wire  [15:0] out_e365;
wire  [15:0] out_e366;
wire  [15:0] out_e367;
wire  [15:0] out_e368;
wire  [15:0] out_e369;
wire  [15:0] out_e370;
wire  [15:0] out_e371;
wire  [15:0] out_e372;
wire  [15:0] out_e373;
wire  [15:0] out_e374;
wire  [15:0] out_e375;
wire  [15:0] out_e376;
wire  [15:0] out_e377;
wire  [15:0] out_e378;
wire  [15:0] out_e379;
wire  [15:0] out_e380;
wire  [15:0] out_e381;
wire  [15:0] out_e382;
wire  [15:0] out_e383;
wire  [15:0] out_e384;
wire  [15:0] out_e385;
wire  [15:0] out_e386;
wire  [15:0] out_e387;
wire  [15:0] out_e388;
wire  [15:0] out_e389;
wire  [15:0] out_e390;
wire  [15:0] out_e391;
wire  [15:0] out_e392;
wire  [15:0] out_e393;
wire  [15:0] out_e394;
wire  [15:0] out_e395;
wire  [15:0] out_e396;
wire  [15:0] out_e397;
wire  [15:0] out_e398;
wire  [15:0] out_e399;
wire  [15:0] out_e400;
wire  [15:0] out_e401;
wire  [15:0] out_e402;
wire  [15:0] out_e403;
wire  [15:0] out_e404;
wire  [15:0] out_e405;
wire  [15:0] out_e406;
wire  [15:0] out_e407;
wire  [15:0] out_e408;
wire  [15:0] out_e409;
wire  [15:0] out_e410;
wire  [15:0] out_e411;
wire  [15:0] out_e412;
wire  [15:0] out_e413;
wire  [15:0] out_e414;
wire  [15:0] out_e415;
wire  [15:0] out_e416;
wire  [15:0] out_e417;
wire  [15:0] out_e418;
wire  [15:0] out_e419;
wire  [15:0] out_e420;
wire  [15:0] out_e421;
wire  [15:0] out_e422;
wire  [15:0] out_e423;
wire  [15:0] out_e424;
wire  [15:0] out_e425;
wire  [15:0] out_e426;
wire  [15:0] out_e427;
wire  [15:0] out_e428;
wire  [15:0] out_e429;
wire  [15:0] out_e430;
wire  [15:0] out_e431;
wire  [15:0] out_e432;
wire  [15:0] out_e433;
wire  [15:0] out_e434;
wire  [15:0] out_e435;
wire  [15:0] out_e436;
wire  [15:0] out_e437;
wire  [15:0] out_e438;
wire  [15:0] out_e439;
wire  [15:0] out_e440;
wire  [15:0] out_e441;
wire  [15:0] out_e442;
wire  [15:0] out_e443;
wire  [15:0] out_e444;
wire  [15:0] out_e445;
wire  [15:0] out_e446;
wire  [15:0] out_e447;
wire  [15:0] out_e448;
wire  [15:0] out_e449;
wire  [15:0] out_e450;
wire  [15:0] out_e451;
wire  [15:0] out_e452;
wire  [15:0] out_e453;
wire  [15:0] out_e454;
wire  [15:0] out_e455;
wire  [15:0] out_e456;
wire  [15:0] out_e457;
wire  [15:0] out_e458;
wire  [15:0] out_e459;
wire  [15:0] out_e460;
wire  [15:0] out_e461;
wire  [15:0] out_e462;
wire  [15:0] out_e463;
wire  [15:0] out_e464;
wire  [15:0] out_e465;
wire  [15:0] out_e466;
wire  [15:0] out_e467;
wire  [15:0] out_e468;
wire  [15:0] out_e469;
wire  [15:0] out_e470;
wire  [15:0] out_e471;
wire  [15:0] out_e472;
wire  [15:0] out_e473;
wire  [15:0] out_e474;
wire  [15:0] out_e475;
wire  [15:0] out_e476;
wire  [15:0] out_e477;
wire  [15:0] out_e478;
wire  [15:0] out_e479;
wire  [15:0] out_e480;
wire  [15:0] out_e481;
wire  [15:0] out_e482;
wire  [15:0] out_e483;
wire  [15:0] out_e484;
wire  [15:0] out_e485;
wire  [15:0] out_e486;
wire  [15:0] out_e487;
wire  [15:0] out_e488;
wire  [15:0] out_e489;
wire  [15:0] out_e490;
wire  [15:0] out_e491;
wire  [15:0] out_e492;
wire  [15:0] out_e493;
wire  [15:0] out_e494;
wire  [15:0] out_e495;
wire  [15:0] out_e496;
wire  [15:0] out_e497;
wire  [15:0] out_e498;
wire  [15:0] out_e499;
wire  [15:0] out_e500;
wire  [15:0] out_e501;
wire  [15:0] out_e502;
wire  [15:0] out_e503;
wire  [15:0] out_e504;
wire  [15:0] out_e505;
wire  [15:0] out_e506;
wire  [15:0] out_e507;
wire  [15:0] out_e508;
wire  [15:0] out_e509;
wire  [15:0] out_e510;
wire  [15:0] out_e511;
wire  [15:0] out_e512;
wire  [15:0] out_e513;
wire  [15:0] out_e514;
wire  [15:0] out_e515;
wire  [15:0] out_e516;
wire  [15:0] out_e517;
wire  [15:0] out_e518;
wire  [15:0] out_e519;
wire  [15:0] out_e520;
wire  [15:0] out_e521;
wire  [15:0] out_e522;
wire  [15:0] out_e523;
wire  [15:0] out_e524;
wire  [15:0] out_e525;
wire  [15:0] out_e526;
wire  [15:0] out_e527;
wire  [15:0] out_e528;
wire  [15:0] out_e529;
wire  [15:0] out_e530;
wire  [15:0] out_e531;
wire  [15:0] out_e532;
wire  [15:0] out_e533;
wire  [15:0] out_e534;
wire  [15:0] out_e535;
wire  [15:0] out_e536;
wire  [15:0] out_e537;
wire  [15:0] out_e538;
wire  [15:0] out_e539;
wire  [15:0] out_e540;
wire  [15:0] out_e541;
wire  [15:0] out_e542;
wire  [15:0] out_e543;
wire  [15:0] out_e544;
wire  [15:0] out_e545;
wire  [15:0] out_e546;
wire  [15:0] out_e547;
wire  [15:0] out_e548;
wire  [15:0] out_e549;
wire  [15:0] out_e550;
wire  [15:0] out_e551;
wire  [15:0] out_e552;
wire  [15:0] out_e553;
wire  [15:0] out_e554;
wire  [15:0] out_e555;
wire  [15:0] out_e556;
wire  [15:0] out_e557;
wire  [15:0] out_e558;
wire  [15:0] out_e559;
wire  [15:0] out_e560;
wire  [15:0] out_e561;
wire  [15:0] out_e562;
wire  [15:0] out_e563;
wire  [15:0] out_e564;
wire  [15:0] out_e565;
wire  [15:0] out_e566;
wire  [15:0] out_e567;
wire  [15:0] out_e568;
wire  [15:0] out_e569;
wire  [15:0] out_e570;
wire  [15:0] out_e571;
wire  [15:0] out_e572;
wire  [15:0] out_e573;
wire  [15:0] out_e574;
wire  [15:0] out_e575;
wire  [15:0] out_e576;
wire  [15:0] out_e577;
wire  [15:0] out_e578;
wire  [15:0] out_e579;
wire  [15:0] out_e580;
wire  [15:0] out_e581;
wire  [15:0] out_e582;
wire  [15:0] out_e583;
wire  [15:0] out_e584;
wire  [15:0] out_e585;
wire  [15:0] out_e586;
wire  [15:0] out_e587;
wire  [15:0] out_e588;
wire  [15:0] out_e589;
wire  [15:0] out_e590;
wire  [15:0] out_e591;
wire  [15:0] out_e592;
wire  [15:0] out_e593;
wire  [15:0] out_e594;
wire  [15:0] out_e595;
wire  [15:0] out_e596;
wire  [15:0] out_e597;
wire  [15:0] out_e598;
wire  [15:0] out_e599;
wire  [15:0] out_e600;
wire  [15:0] out_e601;
wire  [15:0] out_e602;
wire  [15:0] out_e603;
wire  [15:0] out_e604;
wire  [15:0] out_e605;
wire  [15:0] out_e606;
wire  [15:0] out_e607;
wire  [15:0] out_e608;
wire  [15:0] out_e609;
wire  [15:0] out_e610;
wire  [15:0] out_e611;
wire  [15:0] out_e612;
wire  [15:0] out_e613;
wire  [15:0] out_e614;
wire  [15:0] out_e615;
wire  [15:0] out_e616;
wire  [15:0] out_e617;
wire  [15:0] out_e618;
wire  [15:0] out_e619;
wire  [15:0] out_e620;
wire  [15:0] out_e621;
wire  [15:0] out_e622;
wire  [15:0] out_e623;
wire  [15:0] out_e624;
wire  [15:0] out_e625;
wire  [15:0] out_e626;
wire  [15:0] out_e627;
wire  [15:0] out_e628;
wire  [15:0] out_e629;
wire  [15:0] out_e630;
wire  [15:0] out_e631;
wire  [15:0] out_e632;
wire  [15:0] out_e633;
wire  [15:0] out_e634;
wire  [15:0] out_e635;
wire  [15:0] out_e636;
wire  [15:0] out_e637;
wire  [15:0] out_e638;
wire  [15:0] out_e639;
wire  [15:0] out_e640;
wire  [15:0] out_e641;
wire  [15:0] out_e642;
wire  [15:0] out_e643;
wire  [15:0] out_e644;
wire  [15:0] out_e645;
wire  [15:0] out_e646;
wire  [15:0] out_e647;
wire  [15:0] out_e648;
wire  [15:0] out_e649;
wire  [15:0] out_e650;
wire  [15:0] out_e651;
wire  [15:0] out_e652;
wire  [15:0] out_e653;
wire  [15:0] out_e654;
wire  [15:0] out_e655;
wire  [15:0] out_e656;
wire  [15:0] out_e657;
wire  [15:0] out_e658;
wire  [15:0] out_e659;
wire  [15:0] out_e660;
wire  [15:0] out_e661;
wire  [15:0] out_e662;
wire  [15:0] out_e663;
wire  [15:0] out_e664;
wire  [15:0] out_e665;
wire  [15:0] out_e666;
wire  [15:0] out_e667;
wire  [15:0] out_e668;
wire  [15:0] out_e669;
wire  [15:0] out_e670;
wire  [15:0] out_e671;
wire  [15:0] out_e672;
wire  [15:0] out_e673;
wire  [15:0] out_e674;
wire  [15:0] out_e675;
wire  [15:0] out_e676;
wire  [15:0] out_e677;
wire  [15:0] out_e678;
wire  [15:0] out_e679;
wire  [15:0] out_e680;
wire  [15:0] out_e681;
wire  [15:0] out_e682;
wire  [15:0] out_e683;
wire  [15:0] out_e684;
wire  [15:0] out_e685;
wire  [15:0] out_e686;
wire  [15:0] out_e687;
wire  [15:0] out_e688;
wire  [15:0] out_e689;
wire  [15:0] out_e690;
wire  [15:0] out_e691;
wire  [15:0] out_e692;
wire  [15:0] out_e693;
wire  [15:0] out_e694;
wire  [15:0] out_e695;
wire  [15:0] out_e696;
wire  [15:0] out_e697;
wire  [15:0] out_e698;
wire  [15:0] out_e699;
wire  [15:0] out_e700;
wire  [15:0] out_e701;
wire  [15:0] out_e702;
wire  [15:0] out_e703;
wire  [15:0] out_e704;
wire  [15:0] out_e705;
wire  [15:0] out_e706;
wire  [15:0] out_e707;
wire  [15:0] out_e708;
wire  [15:0] out_e709;
wire  [15:0] out_e710;
wire  [15:0] out_e711;
wire  [15:0] out_e712;
wire  [15:0] out_e713;
wire  [15:0] out_e714;
wire  [15:0] out_e715;
wire  [15:0] out_e716;
wire  [15:0] out_e717;
wire  [15:0] out_e718;
wire  [15:0] out_e719;
wire  [15:0] out_e720;
wire  [15:0] out_e721;
wire  [15:0] out_e722;
wire  [15:0] out_e723;
wire  [15:0] out_e724;
wire  [15:0] out_e725;
wire  [15:0] out_e726;
wire  [15:0] out_e727;
wire  [15:0] out_e728;
wire  [15:0] out_e729;
wire  [15:0] out_e730;
wire  [15:0] out_e731;
wire  [15:0] out_e732;
wire  [15:0] out_e733;
wire  [15:0] out_e734;
wire  [15:0] out_e735;
wire  [15:0] out_e736;
wire  [15:0] out_e737;
wire  [15:0] out_e738;
wire  [15:0] out_e739;
wire  [15:0] out_e740;
wire  [15:0] out_e741;
wire  [15:0] out_e742;
wire  [15:0] out_e743;
wire  [15:0] out_e744;
wire  [15:0] out_e745;
wire  [15:0] out_e746;
wire  [15:0] out_e747;
wire  [15:0] out_e748;
wire  [15:0] out_e749;
wire  [15:0] out_e750;
wire  [15:0] out_e751;
wire  [15:0] out_e752;
wire  [15:0] out_e753;
wire  [15:0] out_e754;
wire  [15:0] out_e755;
wire  [15:0] out_e756;
wire  [15:0] out_e757;
wire  [15:0] out_e758;
wire  [15:0] out_e759;
wire  [15:0] out_e760;
wire  [15:0] out_e761;
wire  [15:0] out_e762;
wire  [15:0] out_e763;
wire  [15:0] out_e764;
wire  [15:0] out_e765;
wire  [15:0] out_e766;
wire  [15:0] out_e767;
wire  [15:0] out_e768;
wire  [15:0] out_e769;
wire  [15:0] out_e770;
wire  [15:0] out_e771;
wire  [15:0] out_e772;
wire  [15:0] out_e773;
wire  [15:0] out_e774;
wire  [15:0] out_e775;
wire  [15:0] out_e776;
wire  [15:0] out_e777;
wire  [15:0] out_e778;
wire  [15:0] out_e779;
wire  [15:0] out_e780;
wire  [15:0] out_e781;
wire  [15:0] out_e782;
wire  [15:0] out_e783;
wire  [15:0] out_e784;
wire  [15:0] out_e785;
wire  [15:0] out_e786;
wire  [15:0] out_e787;
wire  [15:0] out_e788;
wire  [15:0] out_e789;
wire  [15:0] out_e790;
wire  [15:0] out_e791;
wire  [15:0] out_e792;
wire  [15:0] out_e793;
wire  [15:0] out_e794;
wire  [15:0] out_e795;
wire  [15:0] out_e796;
wire  [15:0] out_e797;
wire  [15:0] out_e798;
wire  [15:0] out_e799;
wire  [15:0] out_e800;
wire  [15:0] out_e801;
wire  [15:0] out_e802;
wire  [15:0] out_e803;
wire  [15:0] out_e804;
wire  [15:0] out_e805;
wire  [15:0] out_e806;
wire  [15:0] out_e807;
wire  [15:0] out_e808;
wire  [15:0] out_e809;
wire  [15:0] out_e810;
wire  [15:0] out_e811;
wire  [15:0] out_e812;
wire  [15:0] out_e813;
wire  [15:0] out_e814;
wire  [15:0] out_e815;
wire  [15:0] out_e816;
wire  [15:0] out_e817;
wire  [15:0] out_e818;
wire  [15:0] out_e819;
wire  [15:0] out_e820;
wire  [15:0] out_e821;
wire  [15:0] out_e822;
wire  [15:0] out_e823;
wire  [15:0] out_e824;
wire  [15:0] out_e825;
wire  [15:0] out_e826;
wire  [15:0] out_e827;
wire  [15:0] out_e828;
wire  [15:0] out_e829;
wire  [15:0] out_e830;
wire  [15:0] out_e831;
wire  [15:0] out_e832;
wire  [15:0] out_e833;
wire  [15:0] out_e834;
wire  [15:0] out_e835;
wire  [15:0] out_e836;
wire  [15:0] out_e837;
wire  [15:0] out_e838;
wire  [15:0] out_e839;
wire  [15:0] out_e840;
wire  [15:0] out_e841;
wire  [15:0] out_e842;
wire  [15:0] out_e843;
wire  [15:0] out_e844;
wire  [15:0] out_e845;
wire  [15:0] out_e846;
wire  [15:0] out_e847;
wire  [15:0] out_e848;
wire  [15:0] out_e849;
wire  [15:0] out_e850;
wire  [15:0] out_e851;
wire  [15:0] out_e852;
wire  [15:0] out_e853;
wire  [15:0] out_e854;
wire  [15:0] out_e855;
wire  [15:0] out_e856;
wire  [15:0] out_e857;
wire  [15:0] out_e858;
wire  [15:0] out_e859;
wire  [15:0] out_e860;
wire  [15:0] out_e861;
wire  [15:0] out_e862;
wire  [15:0] out_e863;
wire  [15:0] out_e864;
wire  [15:0] out_e865;
wire  [15:0] out_e866;
wire  [15:0] out_e867;
wire  [15:0] out_e868;
wire  [15:0] out_e869;
wire  [15:0] out_e870;
wire  [15:0] out_e871;
wire  [15:0] out_e872;
wire  [15:0] out_e873;
wire  [15:0] out_e874;
wire  [15:0] out_e875;
wire  [15:0] out_e876;
wire  [15:0] out_e877;
wire  [15:0] out_e878;
wire  [15:0] out_e879;
wire  [15:0] out_e880;
wire  [15:0] out_e881;
wire  [15:0] out_e882;
wire  [15:0] out_e883;
wire  [15:0] out_e884;
wire  [15:0] out_e885;
wire  [15:0] out_e886;
wire  [15:0] out_e887;
wire  [15:0] out_e888;
wire  [15:0] out_e889;
wire  [15:0] out_e890;
wire  [15:0] out_e891;
wire  [15:0] out_e892;
wire  [15:0] out_e893;
wire  [15:0] out_e894;
wire  [15:0] out_e895;
wire  [15:0] out_e896;
wire  [15:0] out_e897;
wire  [15:0] out_e898;
wire  [15:0] out_e899;
wire  [15:0] out_e900;
wire  [15:0] out_e901;
wire  [15:0] out_e902;
wire  [15:0] out_e903;
wire  [15:0] out_e904;
wire  [15:0] out_e905;
wire  [15:0] out_e906;
wire  [15:0] out_e907;
wire  [15:0] out_e908;
wire  [15:0] out_e909;
wire  [15:0] out_e910;
wire  [15:0] out_e911;
wire  [15:0] out_e912;
wire  [15:0] out_e913;
wire  [15:0] out_e914;
wire  [15:0] out_e915;
wire  [15:0] out_e916;
wire  [15:0] out_e917;
wire  [15:0] out_e918;
wire  [15:0] out_e919;
wire  [15:0] out_e920;
wire  [15:0] out_e921;
wire  [15:0] out_e922;
wire  [15:0] out_e923;
wire  [15:0] out_e924;
wire  [15:0] out_e925;
wire  [15:0] out_e926;
wire  [15:0] out_e927;
wire  [15:0] out_e928;
wire  [15:0] out_e929;
wire  [15:0] out_e930;
wire  [15:0] out_e931;
wire  [15:0] out_e932;
wire  [15:0] out_e933;
wire  [15:0] out_e934;
wire  [15:0] out_e935;
wire  [15:0] out_e936;
wire  [15:0] out_e937;
wire  [15:0] out_e938;
wire  [15:0] out_e939;
wire  [15:0] out_e940;
wire  [15:0] out_e941;
wire  [15:0] out_e942;
wire  [15:0] out_e943;
wire  [15:0] out_e944;
wire  [15:0] out_e945;
wire  [15:0] out_e946;
wire  [15:0] out_e947;
wire  [15:0] out_e948;
wire  [15:0] out_e949;
wire  [15:0] out_e950;
wire  [15:0] out_e951;
wire  [15:0] out_e952;
wire  [15:0] out_e953;
wire  [15:0] out_e954;
wire  [15:0] out_e955;
wire  [15:0] out_e956;
wire  [15:0] out_e957;
wire  [15:0] out_e958;
wire  [15:0] out_e959;
wire  [15:0] out_e960;
wire  [15:0] out_e961;
wire  [15:0] out_e962;
wire  [15:0] out_e963;
wire  [15:0] out_e964;
wire  [15:0] out_e965;
wire  [15:0] out_e966;
wire  [15:0] out_e967;
wire  [15:0] out_e968;
wire  [15:0] out_e969;
wire  [15:0] out_e970;
wire  [15:0] out_e971;
wire  [15:0] out_e972;
wire  [15:0] out_e973;
wire  [15:0] out_e974;
wire  [15:0] out_e975;
wire  [15:0] out_e976;
wire  [15:0] out_e977;
wire  [15:0] out_e978;
wire  [15:0] out_e979;
wire  [15:0] out_e980;
wire  [15:0] out_e981;
wire  [15:0] out_e982;
wire  [15:0] out_e983;
wire  [15:0] out_e984;
wire  [15:0] out_e985;
wire  [15:0] out_e986;
wire  [15:0] out_e987;
wire  [15:0] out_e988;
wire  [15:0] out_e989;
wire  [15:0] out_e990;
wire  [15:0] out_e991;
wire  [15:0] out_e992;
wire  [15:0] out_e993;
wire  [15:0] out_e994;
wire  [15:0] out_e995;
wire  [15:0] out_e996;
wire  [15:0] out_e997;
wire  [15:0] out_e998;
wire  [15:0] out_e999;
wire  [15:0] out_e1000;
wire  [15:0] out_e1001;
wire  [15:0] out_e1002;
wire  [15:0] out_e1003;
wire  [15:0] out_e1004;
wire  [15:0] out_e1005;
wire  [15:0] out_e1006;
wire  [15:0] out_e1007;
wire  [15:0] out_e1008;
wire  [15:0] out_e1009;
wire  [15:0] out_e1010;
wire  [15:0] out_e1011;
wire  [15:0] out_e1012;
wire  [15:0] out_e1013;
wire  [15:0] out_e1014;
wire  [15:0] out_e1015;
wire  [15:0] out_e1016;
wire  [15:0] out_e1017;
wire  [15:0] out_e1018;
wire  [15:0] out_e1019;
wire  [15:0] out_e1020;
wire  [15:0] out_e1021;
wire  [15:0] out_e1022;
wire  [15:0] out_e1023;
wire  [15:0] out_e1024;
wire  [15:0] out_e1025;
wire  [15:0] out_e1026;
wire  [15:0] out_e1027;
wire  [15:0] out_e1028;
wire  [15:0] out_e1029;
wire  [15:0] out_e1030;
wire  [15:0] out_e1031;
wire  [15:0] out_e1032;
wire  [15:0] out_e1033;
wire  [15:0] out_e1034;
wire  [15:0] out_e1035;
wire  [15:0] out_e1036;
wire  [15:0] out_e1037;
wire  [15:0] out_e1038;
wire  [15:0] out_e1039;
wire  [15:0] out_e1040;
wire  [15:0] out_e1041;
wire  [15:0] out_e1042;
wire  [15:0] out_e1043;
wire  [15:0] out_e1044;
wire  [15:0] out_e1045;
wire  [15:0] out_e1046;
wire  [15:0] out_e1047;
wire  [15:0] out_e1048;
wire  [15:0] out_e1049;
wire  [15:0] out_e1050;
wire  [15:0] out_e1051;
wire  [15:0] out_e1052;
wire  [15:0] out_e1053;
wire  [15:0] out_e1054;
wire  [15:0] out_e1055;
wire  [15:0] out_e1056;
wire  [15:0] out_e1057;
wire  [15:0] out_e1058;
wire  [15:0] out_e1059;
wire  [15:0] out_e1060;
wire  [15:0] out_e1061;
wire  [15:0] out_e1062;
wire  [15:0] out_e1063;
wire  [15:0] out_e1064;
wire  [15:0] out_e1065;
wire  [15:0] out_e1066;
wire  [15:0] out_e1067;
wire  [15:0] out_e1068;
wire  [15:0] out_e1069;
wire  [15:0] out_e1070;
wire  [15:0] out_e1071;
wire  [15:0] out_e1072;
wire  [15:0] out_e1073;
wire  [15:0] out_e1074;
wire  [15:0] out_e1075;
wire  [15:0] out_e1076;
wire  [15:0] out_e1077;
wire  [15:0] out_e1078;
wire  [15:0] out_e1079;
wire  [15:0] out_e1080;
wire  [15:0] out_e1081;
wire  [15:0] out_e1082;
wire  [15:0] out_e1083;
wire  [15:0] out_e1084;
wire  [15:0] out_e1085;
wire  [15:0] out_e1086;
wire  [15:0] out_e1087;
wire  [15:0] out_e1088;
wire  [15:0] out_e1089;
wire  [15:0] out_e1090;
wire  [15:0] out_e1091;
wire  [15:0] out_e1092;
wire  [15:0] out_e1093;
wire  [15:0] out_e1094;
wire  [15:0] out_e1095;
wire  [15:0] out_e1096;
wire  [15:0] out_e1097;
wire  [15:0] out_e1098;
wire  [15:0] out_e1099;
wire  [15:0] out_e1100;
wire  [15:0] out_e1101;
wire  [15:0] out_e1102;
wire  [15:0] out_e1103;
wire  [15:0] out_e1104;
wire  [15:0] out_e1105;
wire  [15:0] out_e1106;
wire  [15:0] out_e1107;
wire  [15:0] out_e1108;
wire  [15:0] out_e1109;
wire  [15:0] out_e1110;
wire  [15:0] out_e1111;
wire  [15:0] out_e1112;
wire  [15:0] out_e1113;
wire  [15:0] out_e1114;
wire  [15:0] out_e1115;
wire  [15:0] out_e1116;
wire  [15:0] out_e1117;
wire  [15:0] out_e1118;
wire  [15:0] out_e1119;
wire  [15:0] out_e1120;
wire  [15:0] out_e1121;
wire  [15:0] out_e1122;
wire  [15:0] out_e1123;
wire  [15:0] out_e1124;
wire  [15:0] out_e1125;
wire  [15:0] out_e1126;
wire  [15:0] out_e1127;
wire  [15:0] out_e1128;
wire  [15:0] out_e1129;
wire  [15:0] out_e1130;
wire  [15:0] out_e1131;
wire  [15:0] out_e1132;
wire  [15:0] out_e1133;
wire  [15:0] out_e1134;
wire  [15:0] out_e1135;
wire  [15:0] out_e1136;
wire  [15:0] out_e1137;
wire  [15:0] out_e1138;
wire  [15:0] out_e1139;
wire  [15:0] out_e1140;
wire  [15:0] out_e1141;
wire  [15:0] out_e1142;
wire  [15:0] out_e1143;
wire  [15:0] out_e1144;
wire  [15:0] out_e1145;
wire  [15:0] out_e1146;
wire  [15:0] out_e1147;
wire  [15:0] out_e1148;
wire  [15:0] out_e1149;
wire  [15:0] out_e1150;
wire  [15:0] out_e1151;
wire  [15:0] out_e1152;
wire  [15:0] out_e1153;
wire  [15:0] out_e1154;
wire  [15:0] out_e1155;
wire  [15:0] out_e1156;
wire  [15:0] out_e1157;
wire  [15:0] out_e1158;
wire  [15:0] out_e1159;
wire  [15:0] out_e1160;
wire  [15:0] out_e1161;
wire  [15:0] out_e1162;
wire  [15:0] out_e1163;
wire  [15:0] out_e1164;
wire  [15:0] out_e1165;
wire  [15:0] out_e1166;
wire  [15:0] out_e1167;
wire  [15:0] out_e1168;
wire  [15:0] out_e1169;
wire  [15:0] out_e1170;
wire  [15:0] out_e1171;
wire  [15:0] out_e1172;
wire  [15:0] out_e1173;
wire  [15:0] out_e1174;
wire  [15:0] out_e1175;
wire  [15:0] out_e1176;
wire  [15:0] out_e1177;
wire  [15:0] out_e1178;
wire  [15:0] out_e1179;
wire  [15:0] out_e1180;
wire  [15:0] out_e1181;
wire  [15:0] out_e1182;
wire  [15:0] out_e1183;
wire  [15:0] out_e1184;
wire  [15:0] out_e1185;
wire  [15:0] out_e1186;
wire  [15:0] out_e1187;
wire  [15:0] out_e1188;
wire  [15:0] out_e1189;
wire  [15:0] out_e1190;
wire  [15:0] out_e1191;
wire  [15:0] out_e1192;
wire  [15:0] out_e1193;
wire  [15:0] out_e1194;
wire  [15:0] out_e1195;
wire  [15:0] out_e1196;
wire  [15:0] out_e1197;
wire  [15:0] out_e1198;
wire  [15:0] out_e1199;
wire  [15:0] out_e1200;
wire  [15:0] out_e1201;
wire  [15:0] out_e1202;
wire  [15:0] out_e1203;
wire  [15:0] out_e1204;
wire  [15:0] out_e1205;
wire  [15:0] out_e1206;
wire  [15:0] out_e1207;
wire  [15:0] out_e1208;
wire  [15:0] out_e1209;
wire  [15:0] out_e1210;
wire  [15:0] out_e1211;
wire  [15:0] out_e1212;
wire  [15:0] out_e1213;
wire  [15:0] out_e1214;
wire  [15:0] out_e1215;
wire  [15:0] out_e1216;
wire  [15:0] out_e1217;
wire  [15:0] out_e1218;
wire  [15:0] out_e1219;
wire  [15:0] out_e1220;
wire  [15:0] out_e1221;
wire  [15:0] out_e1222;
wire  [15:0] out_e1223;
wire  [15:0] out_e1224;
wire  [15:0] out_e1225;
wire  [15:0] out_e1226;
wire  [15:0] out_e1227;
wire  [15:0] out_e1228;
wire  [15:0] out_e1229;
wire  [15:0] out_e1230;
wire  [15:0] out_e1231;
wire  [15:0] out_e1232;
wire  [15:0] out_e1233;
wire  [15:0] out_e1234;
wire  [15:0] out_e1235;
wire  [15:0] out_e1236;
wire  [15:0] out_e1237;
wire  [15:0] out_e1238;
wire  [15:0] out_e1239;
wire  [15:0] out_e1240;
wire  [15:0] out_e1241;
wire  [15:0] out_e1242;
wire  [15:0] out_e1243;
wire  [15:0] out_e1244;
wire  [15:0] out_e1245;
wire  [15:0] out_e1246;
wire  [15:0] out_e1247;
wire  [15:0] out_e1248;
wire  [15:0] out_e1249;
wire  [15:0] out_e1250;
wire  [15:0] out_e1251;
wire  [15:0] out_e1252;
wire  [15:0] out_e1253;
wire  [15:0] out_e1254;
wire  [15:0] out_e1255;
wire  [15:0] out_e1256;
wire  [15:0] out_e1257;
wire  [15:0] out_e1258;
wire  [15:0] out_e1259;
wire  [15:0] out_e1260;
wire  [15:0] out_e1261;
wire  [15:0] out_e1262;
wire  [15:0] out_e1263;
wire  [15:0] out_e1264;
wire  [15:0] out_e1265;
wire  [15:0] out_e1266;
wire  [15:0] out_e1267;
wire  [15:0] out_e1268;
wire  [15:0] out_e1269;
wire  [15:0] out_e1270;
wire  [15:0] out_e1271;
wire  [15:0] out_e1272;
wire  [15:0] out_e1273;
wire  [15:0] out_e1274;
wire  [15:0] out_e1275;
wire  [15:0] out_e1276;
wire  [15:0] out_e1277;
wire  [15:0] out_e1278;
wire  [15:0] out_e1279;
wire  [15:0] out_e1280;
wire  [15:0] out_e1281;
wire  [15:0] out_e1282;
wire  [15:0] out_e1283;
wire  [15:0] out_e1284;
wire  [15:0] out_e1285;
wire  [15:0] out_e1286;
wire  [15:0] out_e1287;
wire  [15:0] out_e1288;
wire  [15:0] out_e1289;
wire  [15:0] out_e1290;
wire  [15:0] out_e1291;
wire  [15:0] out_e1292;
wire  [15:0] out_e1293;
wire  [15:0] out_e1294;
wire  [15:0] out_e1295;
wire  [15:0] out_e1296;
wire  [15:0] out_e1297;
wire  [15:0] out_e1298;
wire  [15:0] out_e1299;
wire  [15:0] out_e1300;
wire  [15:0] out_e1301;
wire  [15:0] out_e1302;
wire  [15:0] out_e1303;
wire  [15:0] out_e1304;
wire  [15:0] out_e1305;
wire  [15:0] out_e1306;
wire  [15:0] out_e1307;
wire  [15:0] out_e1308;
wire  [15:0] out_e1309;
wire  [15:0] out_e1310;
wire  [15:0] out_e1311;
wire  [15:0] out_e1312;
wire  [15:0] out_e1313;
wire  [15:0] out_e1314;
wire  [15:0] out_e1315;
wire  [15:0] out_e1316;
wire  [15:0] out_e1317;
wire  [15:0] out_e1318;
wire  [15:0] out_e1319;
wire  [15:0] out_e1320;
wire  [15:0] out_e1321;
wire  [15:0] out_e1322;
wire  [15:0] out_e1323;
wire  [15:0] out_e1324;
wire  [15:0] out_e1325;
wire  [15:0] out_e1326;
wire  [15:0] out_e1327;
wire  [15:0] out_e1328;
wire  [15:0] out_e1329;
wire  [15:0] out_e1330;
wire  [15:0] out_e1331;
wire  [15:0] out_e1332;
wire  [15:0] out_e1333;
wire  [15:0] out_e1334;
wire  [15:0] out_e1335;
wire  [15:0] out_e1336;
wire  [15:0] out_e1337;
wire  [15:0] out_e1338;
wire  [15:0] out_e1339;
wire  [15:0] out_e1340;
wire  [15:0] out_e1341;
wire  [15:0] out_e1342;
wire  [15:0] out_e1343;
wire  [15:0] out_e1344;
wire  [15:0] out_e1345;
wire  [15:0] out_e1346;
wire  [15:0] out_e1347;
wire  [15:0] out_e1348;
wire  [15:0] out_e1349;
wire  [15:0] out_e1350;
wire  [15:0] out_e1351;
wire  [15:0] out_e1352;
wire  [15:0] out_e1353;
wire  [15:0] out_e1354;
wire  [15:0] out_e1355;
wire  [15:0] out_e1356;
wire  [15:0] out_e1357;
wire  [15:0] out_e1358;
wire  [15:0] out_e1359;
wire  [15:0] out_e1360;
wire  [15:0] out_e1361;
wire  [15:0] out_e1362;
wire  [15:0] out_e1363;
wire  [15:0] out_e1364;
wire  [15:0] out_e1365;
wire  [15:0] out_e1366;
wire  [15:0] out_e1367;
wire  [15:0] out_e1368;
wire  [15:0] out_e1369;
wire  [15:0] out_e1370;
wire  [15:0] out_e1371;
wire  [15:0] out_e1372;
wire  [15:0] out_e1373;
wire  [15:0] out_e1374;
wire  [15:0] out_e1375;
wire  [15:0] out_e1376;
wire  [15:0] out_e1377;
wire  [15:0] out_e1378;
wire  [15:0] out_e1379;
wire  [15:0] out_e1380;
wire  [15:0] out_e1381;
wire  [15:0] out_e1382;
wire  [15:0] out_e1383;
wire  [15:0] out_e1384;
wire  [15:0] out_e1385;
wire  [15:0] out_e1386;
wire  [15:0] out_e1387;
wire  [15:0] out_e1388;
wire  [15:0] out_e1389;
wire  [15:0] out_e1390;
wire  [15:0] out_e1391;
wire  [15:0] out_e1392;
wire  [15:0] out_e1393;
wire  [15:0] out_e1394;
wire  [15:0] out_e1395;
wire  [15:0] out_e1396;
wire  [15:0] out_e1397;
wire  [15:0] out_e1398;
wire  [15:0] out_e1399;
wire  [15:0] out_e1400;
wire  [15:0] out_e1401;
wire  [15:0] out_e1402;
wire  [15:0] out_e1403;
wire  [15:0] out_e1404;
wire  [15:0] out_e1405;
wire  [15:0] out_e1406;
wire  [15:0] out_e1407;
wire  [15:0] out_e1408;
wire  [15:0] out_e1409;
wire  [15:0] out_e1410;
wire  [15:0] out_e1411;
wire  [15:0] out_e1412;
wire  [15:0] out_e1413;
wire  [15:0] out_e1414;
wire  [15:0] out_e1415;
wire  [15:0] out_e1416;
wire  [15:0] out_e1417;
wire  [15:0] out_e1418;
wire  [15:0] out_e1419;
wire  [15:0] out_e1420;
wire  [15:0] out_e1421;
wire  [15:0] out_e1422;
wire  [15:0] out_e1423;
wire  [15:0] out_e1424;
wire  [15:0] out_e1425;
wire  [15:0] out_e1426;
wire  [15:0] out_e1427;
wire  [15:0] out_e1428;
wire  [15:0] out_e1429;
wire  [15:0] out_e1430;
wire  [15:0] out_e1431;
wire  [15:0] out_e1432;
wire  [15:0] out_e1433;
wire  [15:0] out_e1434;
wire  [15:0] out_e1435;
wire  [15:0] out_e1436;
wire  [15:0] out_e1437;
wire  [15:0] out_e1438;
wire  [15:0] out_e1439;
wire  [15:0] out_e1440;
wire  [15:0] out_e1441;
wire  [15:0] out_e1442;
wire  [15:0] out_e1443;
wire  [15:0] out_e1444;
wire  [15:0] out_e1445;
wire  [15:0] out_e1446;
wire  [15:0] out_e1447;
wire  [15:0] out_e1448;
wire  [15:0] out_e1449;
wire  [15:0] out_e1450;
wire  [15:0] out_e1451;
wire  [15:0] out_e1452;
wire  [15:0] out_e1453;
wire  [15:0] out_e1454;
wire  [15:0] out_e1455;
wire  [15:0] out_e1456;
wire  [15:0] out_e1457;
wire  [15:0] out_e1458;
wire  [15:0] out_e1459;
wire  [15:0] out_e1460;
wire  [15:0] out_e1461;
wire  [15:0] out_e1462;
wire  [15:0] out_e1463;
wire  [15:0] out_e1464;
wire  [15:0] out_e1465;
wire  [15:0] out_e1466;
wire  [15:0] out_e1467;
wire  [15:0] out_e1468;
wire  [15:0] out_e1469;
wire  [15:0] out_e1470;
wire  [15:0] out_e1471;
wire  [15:0] out_e1472;
wire  [15:0] out_e1473;
wire  [15:0] out_e1474;
wire  [15:0] out_e1475;
wire  [15:0] out_e1476;
wire  [15:0] out_e1477;
wire  [15:0] out_e1478;
wire  [15:0] out_e1479;
wire  [15:0] out_e1480;
wire  [15:0] out_e1481;
wire  [15:0] out_e1482;
wire  [15:0] out_e1483;
wire  [15:0] out_e1484;
wire  [15:0] out_e1485;
wire  [15:0] out_e1486;
wire  [15:0] out_e1487;
wire  [15:0] out_e1488;
wire  [15:0] out_e1489;
wire  [15:0] out_e1490;
wire  [15:0] out_e1491;
wire  [15:0] out_e1492;
wire  [15:0] out_e1493;
wire  [15:0] out_e1494;
wire  [15:0] out_e1495;
wire  [15:0] out_e1496;
wire  [15:0] out_e1497;
wire  [15:0] out_e1498;
wire  [15:0] out_e1499;
wire  [15:0] out_e1500;
wire  [15:0] out_e1501;
wire  [15:0] out_e1502;
wire  [15:0] out_e1503;
wire  [15:0] out_e1504;
wire  [15:0] out_e1505;
wire  [15:0] out_e1506;
wire  [15:0] out_e1507;
wire  [15:0] out_e1508;
wire  [15:0] out_e1509;
wire  [15:0] out_e1510;
wire  [15:0] out_e1511;
wire  [15:0] out_e1512;
wire  [15:0] out_e1513;
wire  [15:0] out_e1514;
wire  [15:0] out_e1515;
wire  [15:0] out_e1516;
wire  [15:0] out_e1517;
wire  [15:0] out_e1518;
wire  [15:0] out_e1519;
wire  [15:0] out_e1520;
wire  [15:0] out_e1521;
wire  [15:0] out_e1522;
wire  [15:0] out_e1523;
wire  [15:0] out_e1524;
wire  [15:0] out_e1525;
wire  [15:0] out_e1526;
wire  [15:0] out_e1527;
wire  [15:0] out_e1528;
wire  [15:0] out_e1529;
wire  [15:0] out_e1530;
wire  [15:0] out_e1531;
wire  [15:0] out_e1532;
wire  [15:0] out_e1533;
wire  [15:0] out_e1534;
wire  [15:0] out_e1535;
wire  [15:0] out_e1536;
wire  [15:0] out_e1537;
wire  [15:0] out_e1538;
wire  [15:0] out_e1539;
wire  [15:0] out_e1540;
wire  [15:0] out_e1541;
wire  [15:0] out_e1542;
wire  [15:0] out_e1543;
wire  [15:0] out_e1544;
wire  [15:0] out_e1545;
wire  [15:0] out_e1546;
wire  [15:0] out_e1547;
wire  [15:0] out_e1548;
wire  [15:0] out_e1549;
wire  [15:0] out_e1550;
wire  [15:0] out_e1551;
wire  [15:0] out_e1552;
wire  [15:0] out_e1553;
wire  [15:0] out_e1554;
wire  [15:0] out_e1555;
wire  [15:0] out_e1556;
wire  [15:0] out_e1557;
wire  [15:0] out_e1558;
wire  [15:0] out_e1559;
wire  [15:0] out_e1560;
wire  [15:0] out_e1561;
wire  [15:0] out_e1562;
wire  [15:0] out_e1563;
wire  [15:0] out_e1564;
wire  [15:0] out_e1565;
wire  [15:0] out_e1566;
wire  [15:0] out_e1567;
wire  [15:0] out_e1568;
wire  [15:0] out_e1569;
wire  [15:0] out_e1570;
wire  [15:0] out_e1571;
wire  [15:0] out_e1572;
wire  [15:0] out_e1573;
wire  [15:0] out_e1574;
wire  [15:0] out_e1575;
wire  [15:0] out_e1576;
wire  [15:0] out_e1577;
wire  [15:0] out_e1578;
wire  [15:0] out_e1579;
wire  [15:0] out_e1580;
wire  [15:0] out_e1581;
wire  [15:0] out_e1582;
wire  [15:0] out_e1583;
wire  [15:0] out_e1584;
wire  [15:0] out_e1585;
wire  [15:0] out_e1586;
wire  [15:0] out_e1587;
wire  [15:0] out_e1588;
wire  [15:0] out_e1589;
wire  [15:0] out_e1590;
wire  [15:0] out_e1591;
wire  [15:0] out_e1592;
wire  [15:0] out_e1593;
wire  [15:0] out_e1594;
wire  [15:0] out_e1595;
wire  [15:0] out_e1596;
wire  [15:0] out_e1597;
wire  [15:0] out_e1598;
wire  [15:0] out_e1599;
wire  [15:0] out_e1600;
wire  [15:0] out_e1601;
wire  [15:0] out_e1602;
wire  [15:0] out_e1603;
wire  [15:0] out_e1604;
wire  [15:0] out_e1605;
wire  [15:0] out_e1606;
wire  [15:0] out_e1607;
wire  [15:0] out_e1608;
wire  [15:0] out_e1609;
wire  [15:0] out_e1610;
wire  [15:0] out_e1611;
wire  [15:0] out_e1612;
wire  [15:0] out_e1613;
wire  [15:0] out_e1614;
wire  [15:0] out_e1615;
wire  [15:0] out_e1616;
wire  [15:0] out_e1617;
wire  [15:0] out_e1618;
wire  [15:0] out_e1619;
wire  [15:0] out_e1620;
wire  [15:0] out_e1621;
wire  [15:0] out_e1622;
wire  [15:0] out_e1623;
wire  [15:0] out_e1624;
wire  [15:0] out_e1625;
wire  [15:0] out_e1626;
wire  [15:0] out_e1627;
wire  [15:0] out_e1628;
wire  [15:0] out_e1629;
wire  [15:0] out_e1630;
wire  [15:0] out_e1631;
wire  [15:0] out_e1632;
wire  [15:0] out_e1633;
wire  [15:0] out_e1634;
wire  [15:0] out_e1635;
wire  [15:0] out_e1636;
wire  [15:0] out_e1637;
wire  [15:0] out_e1638;
wire  [15:0] out_e1639;
wire  [15:0] out_e1640;
wire  [15:0] out_e1641;
wire  [15:0] out_e1642;
wire  [15:0] out_e1643;
wire  [15:0] out_e1644;
wire  [15:0] out_e1645;
wire  [15:0] out_e1646;
wire  [15:0] out_e1647;
wire  [15:0] out_e1648;
wire  [15:0] out_e1649;
wire  [15:0] out_e1650;
wire  [15:0] out_e1651;
wire  [15:0] out_e1652;
wire  [15:0] out_e1653;
wire  [15:0] out_e1654;
wire  [15:0] out_e1655;
wire  [15:0] out_e1656;
wire  [15:0] out_e1657;
wire  [15:0] out_e1658;
wire  [15:0] out_e1659;
wire  [15:0] out_e1660;
wire  [15:0] out_e1661;
wire  [15:0] out_e1662;
wire  [15:0] out_e1663;
wire  [15:0] out_e1664;
wire  [15:0] out_e1665;
wire  [15:0] out_e1666;
wire  [15:0] out_e1667;
wire  [15:0] out_e1668;
wire  [15:0] out_e1669;
wire  [15:0] out_e1670;
wire  [15:0] out_e1671;
wire  [15:0] out_e1672;
wire  [15:0] out_e1673;
wire  [15:0] out_e1674;
wire  [15:0] out_e1675;
wire  [15:0] out_e1676;
wire  [15:0] out_e1677;
wire  [15:0] out_e1678;
wire  [15:0] out_e1679;
wire  [15:0] out_e1680;
wire  [15:0] out_e1681;
wire  [15:0] out_e1682;
wire  [15:0] out_e1683;
wire  [15:0] out_e1684;
wire  [15:0] out_e1685;
wire  [15:0] out_e1686;
wire  [15:0] out_e1687;
wire  [15:0] out_e1688;
wire  [15:0] out_e1689;
wire  [15:0] out_e1690;
wire  [15:0] out_e1691;
wire  [15:0] out_e1692;
wire  [15:0] out_e1693;
wire  [15:0] out_e1694;
wire  [15:0] out_e1695;
wire  [15:0] out_e1696;
wire  [15:0] out_e1697;
wire  [15:0] out_e1698;
wire  [15:0] out_e1699;
wire  [15:0] out_e1700;
wire  [15:0] out_e1701;
wire  [15:0] out_e1702;
wire  [15:0] out_e1703;
wire  [15:0] out_e1704;
wire  [15:0] out_e1705;
wire  [15:0] out_e1706;
wire  [15:0] out_e1707;
wire  [15:0] out_e1708;
wire  [15:0] out_e1709;
wire  [15:0] out_e1710;
wire  [15:0] out_e1711;
wire  [15:0] out_e1712;
wire  [15:0] out_e1713;
wire  [15:0] out_e1714;
wire  [15:0] out_e1715;
wire  [15:0] out_e1716;
wire  [15:0] out_e1717;
wire  [15:0] out_e1718;
wire  [15:0] out_e1719;
wire  [15:0] out_e1720;
wire  [15:0] out_e1721;
wire  [15:0] out_e1722;
wire  [15:0] out_e1723;
wire  [15:0] out_e1724;
wire  [15:0] out_e1725;
wire  [15:0] out_e1726;
wire  [15:0] out_e1727;
wire  [15:0] out_e1728;
wire  [15:0] out_e1729;
wire  [15:0] out_e1730;
wire  [15:0] out_e1731;
wire  [15:0] out_e1732;
wire  [15:0] out_e1733;
wire  [15:0] out_e1734;
wire  [15:0] out_e1735;
wire  [15:0] out_e1736;
wire  [15:0] out_e1737;
wire  [15:0] out_e1738;
wire  [15:0] out_e1739;
wire  [15:0] out_e1740;
wire  [15:0] out_e1741;
wire  [15:0] out_e1742;
wire  [15:0] out_e1743;
wire  [15:0] out_e1744;
wire  [15:0] out_e1745;
wire  [15:0] out_e1746;
wire  [15:0] out_e1747;
wire  [15:0] out_e1748;
wire  [15:0] out_e1749;
wire  [15:0] out_e1750;
wire  [15:0] out_e1751;
wire  [15:0] out_e1752;
wire  [15:0] out_e1753;
wire  [15:0] out_e1754;
wire  [15:0] out_e1755;
wire  [15:0] out_e1756;
wire  [15:0] out_e1757;
wire  [15:0] out_e1758;
wire  [15:0] out_e1759;
wire  [15:0] out_e1760;
wire  [15:0] out_e1761;
wire  [15:0] out_e1762;
wire  [15:0] out_e1763;
wire  [15:0] out_e1764;
wire  [15:0] out_e1765;
wire  [15:0] out_e1766;
wire  [15:0] out_e1767;
wire  [15:0] out_e1768;
wire  [15:0] out_e1769;
wire  [15:0] out_e1770;
wire  [15:0] out_e1771;
wire  [15:0] out_e1772;
wire  [15:0] out_e1773;
wire  [15:0] out_e1774;
wire  [15:0] out_e1775;
wire  [15:0] out_e1776;
wire  [15:0] out_e1777;
wire  [15:0] out_e1778;
wire  [15:0] out_e1779;
wire  [15:0] out_e1780;
wire  [15:0] out_e1781;
wire  [15:0] out_e1782;
wire  [15:0] out_e1783;
wire  [15:0] out_e1784;
wire  [15:0] out_e1785;
wire  [15:0] out_e1786;
wire  [15:0] out_e1787;
wire  [15:0] out_e1788;
wire  [15:0] out_e1789;
wire  [15:0] out_e1790;
wire  [15:0] out_e1791;
wire  [15:0] out_e1792;
wire  [15:0] out_e1793;
wire  [15:0] out_e1794;
wire  [15:0] out_e1795;
wire  [15:0] out_e1796;
wire  [15:0] out_e1797;
wire  [15:0] out_e1798;
wire  [15:0] out_e1799;
wire  [15:0] out_e1800;
wire  [15:0] out_e1801;
wire  [15:0] out_e1802;
wire  [15:0] out_e1803;
wire  [15:0] out_e1804;
wire  [15:0] out_e1805;
wire  [15:0] out_e1806;
wire  [15:0] out_e1807;
wire  [15:0] out_e1808;
wire  [15:0] out_e1809;
wire  [15:0] out_e1810;
wire  [15:0] out_e1811;
wire  [15:0] out_e1812;
wire  [15:0] out_e1813;
wire  [15:0] out_e1814;
wire  [15:0] out_e1815;
wire  [15:0] out_e1816;
wire  [15:0] out_e1817;
wire  [15:0] out_e1818;
wire  [15:0] out_e1819;
wire  [15:0] out_e1820;
wire  [15:0] out_e1821;
wire  [15:0] out_e1822;
wire  [15:0] out_e1823;
wire  [15:0] out_e1824;
wire  [15:0] out_e1825;
wire  [15:0] out_e1826;
wire  [15:0] out_e1827;
wire  [15:0] out_e1828;
wire  [15:0] out_e1829;
wire  [15:0] out_e1830;
wire  [15:0] out_e1831;
wire  [15:0] out_e1832;
wire  [15:0] out_e1833;
wire  [15:0] out_e1834;
wire  [15:0] out_e1835;
wire  [15:0] out_e1836;
wire  [15:0] out_e1837;
wire  [15:0] out_e1838;
wire  [15:0] out_e1839;
wire  [15:0] out_e1840;
wire  [15:0] out_e1841;
wire  [15:0] out_e1842;
wire  [15:0] out_e1843;
wire  [15:0] out_e1844;
wire  [15:0] out_e1845;
wire  [15:0] out_e1846;
wire  [15:0] out_e1847;
wire  [15:0] out_e1848;
wire  [15:0] out_e1849;
wire  [15:0] out_e1850;
wire  [15:0] out_e1851;
wire  [15:0] out_e1852;
wire  [15:0] out_e1853;
wire  [15:0] out_e1854;
wire  [15:0] out_e1855;
wire  [15:0] out_e1856;
wire  [15:0] out_e1857;
wire  [15:0] out_e1858;
wire  [15:0] out_e1859;
wire  [15:0] out_e1860;
wire  [15:0] out_e1861;
wire  [15:0] out_e1862;
wire  [15:0] out_e1863;
wire  [15:0] out_e1864;
wire  [15:0] out_e1865;
wire  [15:0] out_e1866;
wire  [15:0] out_e1867;
wire  [15:0] out_e1868;
wire  [15:0] out_e1869;
wire  [15:0] out_e1870;
wire  [15:0] out_e1871;
wire  [15:0] out_e1872;
wire  [15:0] out_e1873;
wire  [15:0] out_e1874;
wire  [15:0] out_e1875;
wire  [15:0] out_e1876;
wire  [15:0] out_e1877;
wire  [15:0] out_e1878;
wire  [15:0] out_e1879;
wire  [15:0] out_e1880;
wire  [15:0] out_e1881;
wire  [15:0] out_e1882;
wire  [15:0] out_e1883;
wire  [15:0] out_e1884;
wire  [15:0] out_e1885;
wire  [15:0] out_e1886;
wire  [15:0] out_e1887;
wire  [15:0] out_e1888;
wire  [15:0] out_e1889;
wire  [15:0] out_e1890;
wire  [15:0] out_e1891;
wire  [15:0] out_e1892;
wire  [15:0] out_e1893;
wire  [15:0] out_e1894;
wire  [15:0] out_e1895;
wire  [15:0] out_e1896;
wire  [15:0] out_e1897;
wire  [15:0] out_e1898;
wire  [15:0] out_e1899;
wire  [15:0] out_e1900;
wire  [15:0] out_e1901;
wire  [15:0] out_e1902;
wire  [15:0] out_e1903;
wire  [15:0] out_e1904;
wire  [15:0] out_e1905;
wire  [15:0] out_e1906;
wire  [15:0] out_e1907;
wire  [15:0] out_e1908;
wire  [15:0] out_e1909;
wire  [15:0] out_e1910;
wire  [15:0] out_e1911;
wire  [15:0] out_e1912;
wire  [15:0] out_e1913;
wire  [15:0] out_e1914;
wire  [15:0] out_e1915;
wire  [15:0] out_e1916;
wire  [15:0] out_e1917;
wire  [15:0] out_e1918;
wire  [15:0] out_e1919;
wire  [15:0] out_e1920;
wire  [15:0] out_e1921;
wire  [15:0] out_e1922;
wire  [15:0] out_e1923;
wire  [15:0] out_e1924;
wire  [15:0] out_e1925;
wire  [15:0] out_e1926;
wire  [15:0] out_e1927;
wire  [15:0] out_e1928;
wire  [15:0] out_e1929;
wire  [15:0] out_e1930;
wire  [15:0] out_e1931;
wire  [15:0] out_e1932;
wire  [15:0] out_e1933;
wire  [15:0] out_e1934;
wire  [15:0] out_e1935;
wire  [15:0] out_e1936;
wire  [15:0] out_e1937;
wire  [15:0] out_e1938;
wire  [15:0] out_e1939;
wire  [15:0] out_e1940;
wire  [15:0] out_e1941;
wire  [15:0] out_e1942;
wire  [15:0] out_e1943;
wire  [15:0] out_e1944;
wire  [15:0] out_e1945;
wire  [15:0] out_e1946;
wire  [15:0] out_e1947;
wire  [15:0] out_e1948;
wire  [15:0] out_e1949;
wire  [15:0] out_e1950;
wire  [15:0] out_e1951;
wire  [15:0] out_e1952;
wire  [15:0] out_e1953;
wire  [15:0] out_e1954;
wire  [15:0] out_e1955;
wire  [15:0] out_e1956;
wire  [15:0] out_e1957;
wire  [15:0] out_e1958;
wire  [15:0] out_e1959;
wire  [15:0] out_e1960;
wire  [15:0] out_e1961;
wire  [15:0] out_e1962;
wire  [15:0] out_e1963;
wire  [15:0] out_e1964;
wire  [15:0] out_e1965;
wire  [15:0] out_e1966;
wire  [15:0] out_e1967;
wire  [15:0] out_e1968;
wire  [15:0] out_e1969;
wire  [15:0] out_e1970;
wire  [15:0] out_e1971;
wire  [15:0] out_e1972;
wire  [15:0] out_e1973;
wire  [15:0] out_e1974;
wire  [15:0] out_e1975;
wire  [15:0] out_e1976;
wire  [15:0] out_e1977;
wire  [15:0] out_e1978;
wire  [15:0] out_e1979;
wire  [15:0] out_e1980;
wire  [15:0] out_e1981;
wire  [15:0] out_e1982;
wire  [15:0] out_e1983;
wire  [15:0] out_e1984;
wire  [15:0] out_e1985;
wire  [15:0] out_e1986;
wire  [15:0] out_e1987;
wire  [15:0] out_e1988;
wire  [15:0] out_e1989;
wire  [15:0] out_e1990;
wire  [15:0] out_e1991;
wire  [15:0] out_e1992;
wire  [15:0] out_e1993;
wire  [15:0] out_e1994;
wire  [15:0] out_e1995;
wire  [15:0] out_e1996;
wire  [15:0] out_e1997;
wire  [15:0] out_e1998;
wire  [15:0] out_e1999;
wire  [15:0] out_e2000;
wire  [15:0] out_e2001;
wire  [15:0] out_e2002;
wire  [15:0] out_e2003;
wire  [15:0] out_e2004;
wire  [15:0] out_e2005;
wire  [15:0] out_e2006;
wire  [15:0] out_e2007;
wire  [15:0] out_e2008;
wire  [15:0] out_e2009;
wire  [15:0] out_e2010;
wire  [15:0] out_e2011;
wire  [15:0] out_e2012;
wire  [15:0] out_e2013;
wire  [15:0] out_e2014;
wire  [15:0] out_e2015;
wire  [15:0] out_e2016;
wire  [15:0] out_e2017;
wire  [15:0] out_e2018;
wire  [15:0] out_e2019;
wire  [15:0] out_e2020;
wire  [15:0] out_e2021;
wire  [15:0] out_e2022;
wire  [15:0] out_e2023;
wire  [15:0] out_e2024;
wire  [15:0] out_e2025;
wire  [15:0] out_e2026;
wire  [15:0] out_e2027;
wire  [15:0] out_e2028;
wire  [15:0] out_e2029;
wire  [15:0] out_e2030;
wire  [15:0] out_e2031;
wire  [15:0] out_e2032;
wire  [15:0] out_e2033;
wire  [15:0] out_e2034;
wire  [15:0] out_e2035;
wire  [15:0] out_e2036;
wire  [15:0] out_e2037;
wire  [15:0] out_e2038;
wire  [15:0] out_e2039;
wire  [15:0] out_e2040;
wire  [15:0] out_e2041;
wire  [15:0] out_e2042;
wire  [15:0] out_e2043;
wire  [15:0] out_e2044;
wire  [15:0] out_e2045;
wire  [15:0] out_e2046;
wire  [15:0] out_e2047;
wire  [15:0] out_e2048;
wire  [15:0] out_e2049;
wire  [15:0] out_e2050;
wire  [15:0] out_e2051;
wire  [15:0] out_e2052;
wire  [15:0] out_e2053;
wire  [15:0] out_e2054;
wire  [15:0] out_e2055;
wire  [15:0] out_e2056;
wire  [15:0] out_e2057;
wire  [15:0] out_e2058;
wire  [15:0] out_e2059;
wire  [15:0] out_e2060;
wire  [15:0] out_e2061;
wire  [15:0] out_e2062;
wire  [15:0] out_e2063;
wire  [15:0] out_e2064;
wire  [15:0] out_e2065;
wire  [15:0] out_e2066;
wire  [15:0] out_e2067;
wire  [15:0] out_e2068;
wire  [15:0] out_e2069;
wire  [15:0] out_e2070;
wire  [15:0] out_e2071;
wire  [15:0] out_e2072;
wire  [15:0] out_e2073;
wire  [15:0] out_e2074;
wire  [15:0] out_e2075;
wire  [15:0] out_e2076;
wire  [15:0] out_e2077;
wire  [15:0] out_e2078;
wire  [15:0] out_e2079;
wire  [15:0] out_e2080;
wire  [15:0] out_e2081;
wire  [15:0] out_e2082;
wire  [15:0] out_e2083;
wire  [15:0] out_e2084;
wire  [15:0] out_e2085;
wire  [15:0] out_e2086;
wire  [15:0] out_e2087;
wire  [15:0] out_e2088;
wire  [15:0] out_e2089;
wire  [15:0] out_e2090;
wire  [15:0] out_e2091;
wire  [15:0] out_e2092;
wire  [15:0] out_e2093;
wire  [15:0] out_e2094;
wire  [15:0] out_e2095;
wire  [15:0] out_e2096;
wire  [15:0] out_e2097;
wire  [15:0] out_e2098;
wire  [15:0] out_e2099;
wire  [15:0] out_e2100;
wire  [15:0] out_e2101;
wire  [15:0] out_e2102;
wire  [15:0] out_e2103;
wire  [15:0] out_e2104;
wire  [15:0] out_e2105;
wire  [15:0] out_e2106;
wire  [15:0] out_e2107;
wire  [15:0] out_e2108;
wire  [15:0] out_e2109;
wire  [15:0] out_e2110;
wire  [15:0] out_e2111;
wire  [15:0] out_e2112;
wire  [15:0] out_e2113;
wire  [15:0] out_e2114;
wire  [15:0] out_e2115;
wire  [15:0] out_e2116;
wire  [15:0] out_e2117;
wire  [15:0] out_e2118;
wire  [15:0] out_e2119;
wire  [15:0] out_e2120;
wire  [15:0] out_e2121;
wire  [15:0] out_e2122;
wire  [15:0] out_e2123;
wire  [15:0] out_e2124;
wire  [15:0] out_e2125;
wire  [15:0] out_e2126;
wire  [15:0] out_e2127;
wire  [15:0] out_e2128;
wire  [15:0] out_e2129;
wire  [15:0] out_e2130;
wire  [15:0] out_e2131;
wire  [15:0] out_e2132;
wire  [15:0] out_e2133;
wire  [15:0] out_e2134;
wire  [15:0] out_e2135;
wire  [15:0] out_e2136;
wire  [15:0] out_e2137;
wire  [15:0] out_e2138;
wire  [15:0] out_e2139;
wire  [15:0] out_e2140;
wire  [15:0] out_e2141;
wire  [15:0] out_e2142;
wire  [15:0] out_e2143;
wire  [15:0] out_e2144;
wire  [15:0] out_e2145;
wire  [15:0] out_e2146;
wire  [15:0] out_e2147;
wire  [15:0] out_e2148;
wire  [15:0] out_e2149;
wire  [15:0] out_e2150;
wire  [15:0] out_e2151;
wire  [15:0] out_e2152;
wire  [15:0] out_e2153;
wire  [15:0] out_e2154;
wire  [15:0] out_e2155;
wire  [15:0] out_e2156;
wire  [15:0] out_e2157;
wire  [15:0] out_e2158;
wire  [15:0] out_e2159;
wire  [15:0] out_e2160;
wire  [15:0] out_e2161;
wire  [15:0] out_e2162;
wire  [15:0] out_e2163;
wire  [15:0] out_e2164;
wire  [15:0] out_e2165;
wire  [15:0] out_e2166;
wire  [15:0] out_e2167;
wire  [15:0] out_e2168;
wire  [15:0] out_e2169;
wire  [15:0] out_e2170;
wire  [15:0] out_e2171;
wire  [15:0] out_e2172;
wire  [15:0] out_e2173;
wire  [15:0] out_e2174;
wire  [15:0] out_e2175;
wire  [15:0] out_e2176;
wire  [15:0] out_e2177;
wire  [15:0] out_e2178;
wire  [15:0] out_e2179;
wire  [15:0] out_e2180;
wire  [15:0] out_e2181;
wire  [15:0] out_e2182;
wire  [15:0] out_e2183;
wire  [15:0] out_e2184;
wire  [15:0] out_e2185;
wire  [15:0] out_e2186;
wire  [15:0] out_e2187;
wire  [15:0] out_e2188;
wire  [15:0] out_e2189;
wire  [15:0] out_e2190;
wire  [15:0] out_e2191;
wire  [15:0] out_e2192;
wire  [15:0] out_e2193;
wire  [15:0] out_e2194;
wire  [15:0] out_e2195;
wire  [15:0] out_e2196;
wire  [15:0] out_e2197;
wire  [15:0] out_e2198;
wire  [15:0] out_e2199;
wire  [15:0] out_e2200;
wire  [15:0] out_e2201;
wire  [15:0] out_e2202;
wire  [15:0] out_e2203;
wire  [15:0] out_e2204;
wire  [15:0] out_e2205;
wire  [15:0] out_e2206;
wire  [15:0] out_e2207;
wire  [15:0] out_e2208;
wire  [15:0] out_e2209;
wire  [15:0] out_e2210;
wire  [15:0] out_e2211;
wire  [15:0] out_e2212;
wire  [15:0] out_e2213;
wire  [15:0] out_e2214;
wire  [15:0] out_e2215;
wire  [15:0] out_e2216;
wire  [15:0] out_e2217;
wire  [15:0] out_e2218;
wire  [15:0] out_e2219;
wire  [15:0] out_e2220;
wire  [15:0] out_e2221;
wire  [15:0] out_e2222;
wire  [15:0] out_e2223;
wire  [15:0] out_e2224;
wire  [15:0] out_e2225;
wire  [15:0] out_e2226;
wire  [15:0] out_e2227;
wire  [15:0] out_e2228;
wire  [15:0] out_e2229;
wire  [15:0] out_e2230;
wire  [15:0] out_e2231;
wire  [15:0] out_e2232;
wire  [15:0] out_e2233;
wire  [15:0] out_e2234;
wire  [15:0] out_e2235;
wire  [15:0] out_e2236;
wire  [15:0] out_e2237;
wire  [15:0] out_e2238;
wire  [15:0] out_e2239;
wire  [15:0] out_e2240;
wire  [15:0] out_e2241;
wire  [15:0] out_e2242;
wire  [15:0] out_e2243;
wire  [15:0] out_e2244;
wire  [15:0] out_e2245;
wire  [15:0] out_e2246;
wire  [15:0] out_e2247;
wire  [15:0] out_e2248;
wire  [15:0] out_e2249;
wire  [15:0] out_e2250;
wire  [15:0] out_e2251;
wire  [15:0] out_e2252;
wire  [15:0] out_e2253;
wire  [15:0] out_e2254;
wire  [15:0] out_e2255;
wire  [15:0] out_e2256;
wire  [15:0] out_e2257;
wire  [15:0] out_e2258;
wire  [15:0] out_e2259;
wire  [15:0] out_e2260;
wire  [15:0] out_e2261;
wire  [15:0] out_e2262;
wire  [15:0] out_e2263;
wire  [15:0] out_e2264;
wire  [15:0] out_e2265;
wire  [15:0] out_e2266;
wire  [15:0] out_e2267;
wire  [15:0] out_e2268;
wire  [15:0] out_e2269;
wire  [15:0] out_e2270;
wire  [15:0] out_e2271;
wire  [15:0] out_e2272;
wire  [15:0] out_e2273;
wire  [15:0] out_e2274;
wire  [15:0] out_e2275;
wire  [15:0] out_e2276;
wire  [15:0] out_e2277;
wire  [15:0] out_e2278;
wire  [15:0] out_e2279;
wire  [15:0] out_e2280;
wire  [15:0] out_e2281;
wire  [15:0] out_e2282;
wire  [15:0] out_e2283;
wire  [15:0] out_e2284;
wire  [15:0] out_e2285;
wire  [15:0] out_e2286;
wire  [15:0] out_e2287;
wire  [15:0] out_e2288;
wire  [15:0] out_e2289;
wire  [15:0] out_e2290;
wire  [15:0] out_e2291;
wire  [15:0] out_e2292;
wire  [15:0] out_e2293;
wire  [15:0] out_e2294;
wire  [15:0] out_e2295;
wire  [15:0] out_e2296;
wire  [15:0] out_e2297;
wire  [15:0] out_e2298;
wire  [15:0] out_e2299;
wire  [15:0] out_e2300;
wire  [15:0] out_e2301;
wire  [15:0] out_e2302;
wire  [15:0] out_e2303;
wire  [15:0] out_e2304;
wire  [15:0] out_e2305;
wire  [15:0] out_e2306;
wire  [15:0] out_e2307;
wire  [15:0] out_e2308;
wire  [15:0] out_e2309;
wire  [15:0] out_e2310;
wire  [15:0] out_e2311;
wire  [15:0] out_e2312;
wire  [15:0] out_e2313;
wire  [15:0] out_e2314;
wire  [15:0] out_e2315;
wire  [15:0] out_e2316;
wire  [15:0] out_e2317;
wire  [15:0] out_e2318;
wire  [15:0] out_e2319;
wire  [15:0] out_e2320;
wire  [15:0] out_e2321;
wire  [15:0] out_e2322;
wire  [15:0] out_e2323;
wire  [15:0] out_e2324;
wire  [15:0] out_e2325;
wire  [15:0] out_e2326;
wire  [15:0] out_e2327;
wire  [15:0] out_e2328;
wire  [15:0] out_e2329;
wire  [15:0] out_e2330;
wire  [15:0] out_e2331;
wire  [15:0] out_e2332;
wire  [15:0] out_e2333;
wire  [15:0] out_e2334;
wire  [15:0] out_e2335;
wire  [15:0] out_e2336;
wire  [15:0] out_e2337;
wire  [15:0] out_e2338;
wire  [15:0] out_e2339;
wire  [15:0] out_e2340;
wire  [15:0] out_e2341;
wire  [15:0] out_e2342;
wire  [15:0] out_e2343;
wire  [15:0] out_e2344;
wire  [15:0] out_e2345;
wire  [15:0] out_e2346;
wire  [15:0] out_e2347;
wire  [15:0] out_e2348;
wire  [15:0] out_e2349;
wire  [15:0] out_e2350;
wire  [15:0] out_e2351;
wire  [15:0] out_e2352;
wire  [15:0] out_e2353;
wire  [15:0] out_e2354;
wire  [15:0] out_e2355;
wire  [15:0] out_e2356;
wire  [15:0] out_e2357;
wire  [15:0] out_e2358;
wire  [15:0] out_e2359;
wire  [15:0] out_e2360;
wire  [15:0] out_e2361;
wire  [15:0] out_e2362;
wire  [15:0] out_e2363;
wire  [15:0] out_e2364;
wire  [15:0] out_e2365;
wire  [15:0] out_e2366;
wire  [15:0] out_e2367;
wire  [15:0] out_e2368;
wire  [15:0] out_e2369;
wire  [15:0] out_e2370;
wire  [15:0] out_e2371;
wire  [15:0] out_e2372;
wire  [15:0] out_e2373;
wire  [15:0] out_e2374;
wire  [15:0] out_e2375;
wire  [15:0] out_e2376;
wire  [15:0] out_e2377;
wire  [15:0] out_e2378;
wire  [15:0] out_e2379;
wire  [15:0] out_e2380;
wire  [15:0] out_e2381;
wire  [15:0] out_e2382;
wire  [15:0] out_e2383;
wire  [15:0] out_e2384;
wire  [15:0] out_e2385;
wire  [15:0] out_e2386;
wire  [15:0] out_e2387;
wire  [15:0] out_e2388;
wire  [15:0] out_e2389;
wire  [15:0] out_e2390;
wire  [15:0] out_e2391;
wire  [15:0] out_e2392;
wire  [15:0] out_e2393;
wire  [15:0] out_e2394;
wire  [15:0] out_e2395;
wire  [15:0] out_e2396;
wire  [15:0] out_e2397;
wire  [15:0] out_e2398;
wire  [15:0] out_e2399;
wire  [15:0] out_e2400;
wire  [15:0] out_e2401;
wire  [15:0] out_e2402;
wire  [15:0] out_e2403;
wire  [15:0] out_e2404;
wire  [15:0] out_e2405;
wire  [15:0] out_e2406;
wire  [15:0] out_e2407;
wire  [15:0] out_e2408;
wire  [15:0] out_e2409;
wire  [15:0] out_e2410;
wire  [15:0] out_e2411;
wire  [15:0] out_e2412;
wire  [15:0] out_e2413;
wire  [15:0] out_e2414;
wire  [15:0] out_e2415;
wire  [15:0] out_e2416;
wire  [15:0] out_e2417;
wire  [15:0] out_e2418;
wire  [15:0] out_e2419;
wire  [15:0] out_e2420;
wire  [15:0] out_e2421;
wire  [15:0] out_e2422;
wire  [15:0] out_e2423;
wire  [15:0] out_e2424;
wire  [15:0] out_e2425;
wire  [15:0] out_e2426;
wire  [15:0] out_e2427;
wire  [15:0] out_e2428;
wire  [15:0] out_e2429;
wire  [15:0] out_e2430;
wire  [15:0] out_e2431;
wire  [15:0] out_e2432;
wire  [15:0] out_e2433;
wire  [15:0] out_e2434;
wire  [15:0] out_e2435;
wire  [15:0] out_e2436;
wire  [15:0] out_e2437;
wire  [15:0] out_e2438;
wire  [15:0] out_e2439;
wire  [15:0] out_e2440;
wire  [15:0] out_e2441;
wire  [15:0] out_e2442;
wire  [15:0] out_e2443;
wire  [15:0] out_e2444;
wire  [15:0] out_e2445;
wire  [15:0] out_e2446;
wire  [15:0] out_e2447;
wire  [15:0] out_e2448;
wire  [15:0] out_e2449;
wire  [15:0] out_e2450;
wire  [15:0] out_e2451;
wire  [15:0] out_e2452;
wire  [15:0] out_e2453;
wire  [15:0] out_e2454;
wire  [15:0] out_e2455;
wire  [15:0] out_e2456;
wire  [15:0] out_e2457;
wire  [15:0] out_e2458;
wire  [15:0] out_e2459;
wire  [15:0] out_e2460;
wire  [15:0] out_e2461;
wire  [15:0] out_e2462;
wire  [15:0] out_e2463;
wire  [15:0] out_e2464;
wire  [15:0] out_e2465;
wire  [15:0] out_e2466;
wire  [15:0] out_e2467;
wire  [15:0] out_e2468;
wire  [15:0] out_e2469;
wire  [15:0] out_e2470;
wire  [15:0] out_e2471;
wire  [15:0] out_e2472;
wire  [15:0] out_e2473;
wire  [15:0] out_e2474;
wire  [15:0] out_e2475;
wire  [15:0] out_e2476;
wire  [15:0] out_e2477;
wire  [15:0] out_e2478;
wire  [15:0] out_e2479;
wire  [15:0] out_e2480;
wire  [15:0] out_e2481;
wire  [15:0] out_e2482;
wire  [15:0] out_e2483;
wire  [15:0] out_e2484;
wire  [15:0] out_e2485;
wire  [15:0] out_e2486;
wire  [15:0] out_e2487;
wire  [15:0] out_e2488;
wire  [15:0] out_e2489;
wire  [15:0] out_e2490;
wire  [15:0] out_e2491;
wire  [15:0] out_e2492;
wire  [15:0] out_e2493;
wire  [15:0] out_e2494;
wire  [15:0] out_e2495;
wire  [15:0] out_e2496;
wire  [15:0] out_e2497;
wire  [15:0] out_e2498;
wire  [15:0] out_e2499;
wire  [15:0] out_e2500;
wire  [15:0] out_e2501;
wire  [15:0] out_e2502;
wire  [15:0] out_e2503;
wire  [15:0] out_e2504;
wire  [15:0] out_e2505;
wire  [15:0] out_e2506;
wire  [15:0] out_e2507;
wire  [15:0] out_e2508;
wire  [15:0] out_e2509;
wire  [15:0] out_e2510;
wire  [15:0] out_e2511;
wire  [15:0] out_e2512;
wire  [15:0] out_e2513;
wire  [15:0] out_e2514;
wire  [15:0] out_e2515;
wire  [15:0] out_e2516;
wire  [15:0] out_e2517;
wire  [15:0] out_e2518;
wire  [15:0] out_e2519;
wire  [15:0] out_e2520;
wire  [15:0] out_e2521;
wire  [15:0] out_e2522;
wire  [15:0] out_e2523;
wire  [15:0] out_e2524;
wire  [15:0] out_e2525;
wire  [15:0] out_e2526;
wire  [15:0] out_e2527;
wire  [15:0] out_e2528;
wire  [15:0] out_e2529;
wire  [15:0] out_e2530;
wire  [15:0] out_e2531;
wire  [15:0] out_e2532;
wire  [15:0] out_e2533;
wire  [15:0] out_e2534;
wire  [15:0] out_e2535;
wire  [15:0] out_e2536;
wire  [15:0] out_e2537;
wire  [15:0] out_e2538;
wire  [15:0] out_e2539;
wire  [15:0] out_e2540;
wire  [15:0] out_e2541;
wire  [15:0] out_e2542;
wire  [15:0] out_e2543;
wire  [15:0] out_e2544;
wire  [15:0] out_e2545;
wire  [15:0] out_e2546;
wire  [15:0] out_e2547;
wire  [15:0] out_e2548;
wire  [15:0] out_e2549;
wire  [15:0] out_e2550;
wire  [15:0] out_e2551;
wire  [15:0] out_e2552;
wire  [15:0] out_e2553;
wire  [15:0] out_e2554;
wire  [15:0] out_e2555;
wire  [15:0] out_e2556;
wire  [15:0] out_e2557;
wire  [15:0] out_e2558;
wire  [15:0] out_e2559;
wire  [15:0] out_e2560;
wire  [15:0] out_e2561;
wire  [15:0] out_e2562;
wire  [15:0] out_e2563;
wire  [15:0] out_e2564;
wire  [15:0] out_e2565;
wire  [15:0] out_e2566;
wire  [15:0] out_e2567;
wire  [15:0] out_e2568;
wire  [15:0] out_e2569;
wire  [15:0] out_e2570;
wire  [15:0] out_e2571;
wire  [15:0] out_e2572;
wire  [15:0] out_e2573;
wire  [15:0] out_e2574;
wire  [15:0] out_e2575;
wire  [15:0] out_e2576;
wire  [15:0] out_e2577;
wire  [15:0] out_e2578;
wire  [15:0] out_e2579;
wire  [15:0] out_e2580;
wire  [15:0] out_e2581;
wire  [15:0] out_e2582;
wire  [15:0] out_e2583;
wire  [15:0] out_e2584;
wire  [15:0] out_e2585;
wire  [15:0] out_e2586;
wire  [15:0] out_e2587;
wire  [15:0] out_e2588;
wire  [15:0] out_e2589;
wire  [15:0] out_e2590;
wire  [15:0] out_e2591;
wire  [15:0] out_e2592;
wire  [15:0] out_e2593;
wire  [15:0] out_e2594;
wire  [15:0] out_e2595;
wire  [15:0] out_e2596;
wire  [15:0] out_e2597;
wire  [15:0] out_e2598;
wire  [15:0] out_e2599;
wire  [15:0] out_e2600;
wire  [15:0] out_e2601;
wire  [15:0] out_e2602;
wire  [15:0] out_e2603;
wire  [15:0] out_e2604;
wire  [15:0] out_e2605;
wire  [15:0] out_e2606;
wire  [15:0] out_e2607;
wire  [15:0] out_e2608;
wire  [15:0] out_e2609;
wire  [15:0] out_e2610;
wire  [15:0] out_e2611;
wire  [15:0] out_e2612;
wire  [15:0] out_e2613;
wire  [15:0] out_e2614;
wire  [15:0] out_e2615;
wire  [15:0] out_e2616;
wire  [15:0] out_e2617;
wire  [15:0] out_e2618;
wire  [15:0] out_e2619;
wire  [15:0] out_e2620;
wire  [15:0] out_e2621;
wire  [15:0] out_e2622;
wire  [15:0] out_e2623;
wire  [15:0] out_e2624;
wire  [15:0] out_e2625;
wire  [15:0] out_e2626;
wire  [15:0] out_e2627;
wire  [15:0] out_e2628;
wire  [15:0] out_e2629;
wire  [15:0] out_e2630;
wire  [15:0] out_e2631;
wire  [15:0] out_e2632;
wire  [15:0] out_e2633;
wire  [15:0] out_e2634;
wire  [15:0] out_e2635;
wire  [15:0] out_e2636;
wire  [15:0] out_e2637;
wire  [15:0] out_e2638;
wire  [15:0] out_e2639;
wire  [15:0] out_e2640;
wire  [15:0] out_e2641;
wire  [15:0] out_e2642;
wire  [15:0] out_e2643;
wire  [15:0] out_e2644;
wire  [15:0] out_e2645;
wire  [15:0] out_e2646;
wire  [15:0] out_e2647;
wire  [15:0] out_e2648;
wire  [15:0] out_e2649;
wire  [15:0] out_e2650;
wire  [15:0] out_e2651;
wire  [15:0] out_e2652;
wire  [15:0] out_e2653;
wire  [15:0] out_e2654;
wire  [15:0] out_e2655;
wire  [15:0] out_e2656;
wire  [15:0] out_e2657;
wire  [15:0] out_e2658;
wire  [15:0] out_e2659;
wire  [15:0] out_e2660;
wire  [15:0] out_e2661;
wire  [15:0] out_e2662;
wire  [15:0] out_e2663;
wire  [15:0] out_e2664;
wire  [15:0] out_e2665;
wire  [15:0] out_e2666;
wire  [15:0] out_e2667;
wire  [15:0] out_e2668;
wire  [15:0] out_e2669;
wire  [15:0] out_e2670;
wire  [15:0] out_e2671;
wire  [15:0] out_e2672;
wire  [15:0] out_e2673;
wire  [15:0] out_e2674;
wire  [15:0] out_e2675;
wire  [15:0] out_e2676;
wire  [15:0] out_e2677;
wire  [15:0] out_e2678;
wire  [15:0] out_e2679;
wire  [15:0] out_e2680;
wire  [15:0] out_e2681;
wire  [15:0] out_e2682;
wire  [15:0] out_e2683;
wire  [15:0] out_e2684;
wire  [15:0] out_e2685;
wire  [15:0] out_e2686;
wire  [15:0] out_e2687;
wire  [15:0] out_e2688;
wire  [15:0] out_e2689;
wire  [15:0] out_e2690;
wire  [15:0] out_e2691;
wire  [15:0] out_e2692;
wire  [15:0] out_e2693;
wire  [15:0] out_e2694;
wire  [15:0] out_e2695;
wire  [15:0] out_e2696;
wire  [15:0] out_e2697;
wire  [15:0] out_e2698;
wire  [15:0] out_e2699;
wire  [15:0] out_e2700;
wire  [15:0] out_e2701;
wire  [15:0] out_e2702;
wire  [15:0] out_e2703;
wire  [15:0] out_e2704;
wire  [15:0] out_e2705;
wire  [15:0] out_e2706;
wire  [15:0] out_e2707;
wire  [15:0] out_e2708;
wire  [15:0] out_e2709;
wire  [15:0] out_e2710;
wire  [15:0] out_e2711;
wire  [15:0] out_e2712;
wire  [15:0] out_e2713;
wire  [15:0] out_e2714;
wire  [15:0] out_e2715;
wire  [15:0] out_e2716;
wire  [15:0] out_e2717;
wire  [15:0] out_e2718;
wire  [15:0] out_e2719;
wire  [15:0] out_e2720;
wire  [15:0] out_e2721;
wire  [15:0] out_e2722;
wire  [15:0] out_e2723;
wire  [15:0] out_e2724;
wire  [15:0] out_e2725;
wire  [15:0] out_e2726;
wire  [15:0] out_e2727;
wire  [15:0] out_e2728;
wire  [15:0] out_e2729;
wire  [15:0] out_e2730;
wire  [15:0] out_e2731;
wire  [15:0] out_e2732;
wire  [15:0] out_e2733;
wire  [15:0] out_e2734;
wire  [15:0] out_e2735;
wire  [15:0] out_e2736;
wire  [15:0] out_e2737;
wire  [15:0] out_e2738;
wire  [15:0] out_e2739;
wire  [15:0] out_e2740;
wire  [15:0] out_e2741;
wire  [15:0] out_e2742;
wire  [15:0] out_e2743;
wire  [15:0] out_e2744;
wire  [15:0] out_e2745;
wire  [15:0] out_e2746;
wire  [15:0] out_e2747;
wire  [15:0] out_e2748;
wire  [15:0] out_e2749;
wire  [15:0] out_e2750;
wire  [15:0] out_e2751;
wire  [15:0] out_e2752;
wire  [15:0] out_e2753;
wire  [15:0] out_e2754;
wire  [15:0] out_e2755;
wire  [15:0] out_e2756;
wire  [15:0] out_e2757;
wire  [15:0] out_e2758;
wire  [15:0] out_e2759;
wire  [15:0] out_e2760;
wire  [15:0] out_e2761;
wire  [15:0] out_e2762;
wire  [15:0] out_e2763;
wire  [15:0] out_e2764;
wire  [15:0] out_e2765;
wire  [15:0] out_e2766;
wire  [15:0] out_e2767;
wire  [15:0] out_e2768;
wire  [15:0] out_e2769;
wire  [15:0] out_e2770;
wire  [15:0] out_e2771;
wire  [15:0] out_e2772;
wire  [15:0] out_e2773;
wire  [15:0] out_e2774;
wire  [15:0] out_e2775;
wire  [15:0] out_e2776;
wire  [15:0] out_e2777;
wire  [15:0] out_e2778;
wire  [15:0] out_e2779;
wire  [15:0] out_e2780;
wire  [15:0] out_e2781;
wire  [15:0] out_e2782;
wire  [15:0] out_e2783;
wire  [15:0] out_e2784;
wire  [15:0] out_e2785;
wire  [15:0] out_e2786;
wire  [15:0] out_e2787;
wire  [15:0] out_e2788;
wire  [15:0] out_e2789;
wire  [15:0] out_e2790;
wire  [15:0] out_e2791;
wire  [15:0] out_e2792;
wire  [15:0] out_e2793;
wire  [15:0] out_e2794;
wire  [15:0] out_e2795;
wire  [15:0] out_e2796;
wire  [15:0] out_e2797;
wire  [15:0] out_e2798;
wire  [15:0] out_e2799;
wire  [15:0] out_e2800;
wire  [15:0] out_e2801;
wire  [15:0] out_e2802;
wire  [15:0] out_e2803;
wire  [15:0] out_e2804;
wire  [15:0] out_e2805;
wire  [15:0] out_e2806;
wire  [15:0] out_e2807;
wire  [15:0] out_e2808;
wire  [15:0] out_e2809;
wire  [15:0] out_e2810;
wire  [15:0] out_e2811;
wire  [15:0] out_e2812;
wire  [15:0] out_e2813;
wire  [15:0] out_e2814;
wire  [15:0] out_e2815;
wire  [15:0] out_e2816;
wire  [15:0] out_e2817;
wire  [15:0] out_e2818;
wire  [15:0] out_e2819;
wire  [15:0] out_e2820;
wire  [15:0] out_e2821;
wire  [15:0] out_e2822;
wire  [15:0] out_e2823;
wire  [15:0] out_e2824;
wire  [15:0] out_e2825;
wire  [15:0] out_e2826;
wire  [15:0] out_e2827;
wire  [15:0] out_e2828;
wire  [15:0] out_e2829;
wire  [15:0] out_e2830;
wire  [15:0] out_e2831;
wire  [15:0] out_e2832;
wire  [15:0] out_e2833;
wire  [15:0] out_e2834;
wire  [15:0] out_e2835;
wire  [15:0] out_e2836;
wire  [15:0] out_e2837;
wire  [15:0] out_e2838;
wire  [15:0] out_e2839;
wire  [15:0] out_e2840;
wire  [15:0] out_e2841;
wire  [15:0] out_e2842;
wire  [15:0] out_e2843;
wire  [15:0] out_e2844;
wire  [15:0] out_e2845;
wire  [15:0] out_e2846;
wire  [15:0] out_e2847;
wire  [15:0] out_e2848;
wire  [15:0] out_e2849;
wire  [15:0] out_e2850;
wire  [15:0] out_e2851;
wire  [15:0] out_e2852;
wire  [15:0] out_e2853;
wire  [15:0] out_e2854;
wire  [15:0] out_e2855;
wire  [15:0] out_e2856;
wire  [15:0] out_e2857;
wire  [15:0] out_e2858;
wire  [15:0] out_e2859;
wire  [15:0] out_e2860;
wire  [15:0] out_e2861;
wire  [15:0] out_e2862;
wire  [15:0] out_e2863;
wire  [15:0] out_e2864;
wire  [15:0] out_e2865;
wire  [15:0] out_e2866;
wire  [15:0] out_e2867;
wire  [15:0] out_e2868;
wire  [15:0] out_e2869;
wire  [15:0] out_e2870;
wire  [15:0] out_e2871;
wire  [15:0] out_e2872;
wire  [15:0] out_e2873;
wire  [15:0] out_e2874;
wire  [15:0] out_e2875;
wire  [15:0] out_e2876;
wire  [15:0] out_e2877;
wire  [15:0] out_e2878;
wire  [15:0] out_e2879;
wire  [15:0] out_e2880;
wire  [15:0] out_e2881;
wire  [15:0] out_e2882;
wire  [15:0] out_e2883;
wire  [15:0] out_e2884;
wire  [15:0] out_e2885;
wire  [15:0] out_e2886;
wire  [15:0] out_e2887;
wire  [15:0] out_e2888;
wire  [15:0] out_e2889;
wire  [15:0] out_e2890;
wire  [15:0] out_e2891;
wire  [15:0] out_e2892;
wire  [15:0] out_e2893;
wire  [15:0] out_e2894;
wire  [15:0] out_e2895;
wire  [15:0] out_e2896;
wire  [15:0] out_e2897;
wire  [15:0] out_e2898;
wire  [15:0] out_e2899;
wire  [15:0] out_e2900;
wire  [15:0] out_e2901;
wire  [15:0] out_e2902;
wire  [15:0] out_e2903;
wire  [15:0] out_e2904;
wire  [15:0] out_e2905;
wire  [15:0] out_e2906;
wire  [15:0] out_e2907;
wire  [15:0] out_e2908;
wire  [15:0] out_e2909;
wire  [15:0] out_e2910;
wire  [15:0] out_e2911;
wire  [15:0] out_e2912;
wire  [15:0] out_e2913;
wire  [15:0] out_e2914;
wire  [15:0] out_e2915;
wire  [15:0] out_e2916;
wire  [15:0] out_e2917;
wire  [15:0] out_e2918;
wire  [15:0] out_e2919;
wire  [15:0] out_e2920;
wire  [15:0] out_e2921;
wire  [15:0] out_e2922;
wire  [15:0] out_e2923;
wire  [15:0] out_e2924;
wire  [15:0] out_e2925;
wire  [15:0] out_e2926;
wire  [15:0] out_e2927;
wire  [15:0] out_e2928;
wire  [15:0] out_e2929;
wire  [15:0] out_e2930;
wire  [15:0] out_e2931;
wire  [15:0] out_e2932;
wire  [15:0] out_e2933;
wire  [15:0] out_e2934;
wire  [15:0] out_e2935;
wire  [15:0] out_e2936;
wire  [15:0] out_e2937;
wire  [15:0] out_e2938;
wire  [15:0] out_e2939;
wire  [15:0] out_e2940;
wire  [15:0] out_e2941;
wire  [15:0] out_e2942;
wire  [15:0] out_e2943;
wire  [15:0] out_e2944;
wire  [15:0] out_e2945;
wire  [15:0] out_e2946;
wire  [15:0] out_e2947;
wire  [15:0] out_e2948;
wire  [15:0] out_e2949;
wire  [15:0] out_e2950;
wire  [15:0] out_e2951;
wire  [15:0] out_e2952;
wire  [15:0] out_e2953;
wire  [15:0] out_e2954;
wire  [15:0] out_e2955;
wire  [15:0] out_e2956;
wire  [15:0] out_e2957;
wire  [15:0] out_e2958;
wire  [15:0] out_e2959;
wire  [15:0] out_e2960;
wire  [15:0] out_e2961;
wire  [15:0] out_e2962;
wire  [15:0] out_e2963;
wire  [15:0] out_e2964;
wire  [15:0] out_e2965;
wire  [15:0] out_e2966;
wire  [15:0] out_e2967;
wire  [15:0] out_e2968;
wire  [15:0] out_e2969;
wire  [15:0] out_e2970;
wire  [15:0] out_e2971;
wire  [15:0] out_e2972;
wire  [15:0] out_e2973;
wire  [15:0] out_e2974;
wire  [15:0] out_e2975;
wire  [15:0] out_e2976;
wire  [15:0] out_e2977;
wire  [15:0] out_e2978;
wire  [15:0] out_e2979;
wire  [15:0] out_e2980;
wire  [15:0] out_e2981;
wire  [15:0] out_e2982;
wire  [15:0] out_e2983;
wire  [15:0] out_e2984;
wire  [15:0] out_e2985;
wire  [15:0] out_e2986;
wire  [15:0] out_e2987;
wire  [15:0] out_e2988;
wire  [15:0] out_e2989;
wire  [15:0] out_e2990;
wire  [15:0] out_e2991;
wire  [15:0] out_e2992;
wire  [15:0] out_e2993;
wire  [15:0] out_e2994;
wire  [15:0] out_e2995;
wire  [15:0] out_e2996;
wire  [15:0] out_e2997;
wire  [15:0] out_e2998;
wire  [15:0] out_e2999;
wire  [15:0] out_e3000;
wire  [15:0] out_e3001;
wire  [15:0] out_e3002;
wire  [15:0] out_e3003;
wire  [15:0] out_e3004;
wire  [15:0] out_e3005;
wire  [15:0] out_e3006;
wire  [15:0] out_e3007;
wire  [15:0] out_e3008;
wire  [15:0] out_e3009;
wire  [15:0] out_e3010;
wire  [15:0] out_e3011;
wire  [15:0] out_e3012;
wire  [15:0] out_e3013;
wire  [15:0] out_e3014;
wire  [15:0] out_e3015;
wire  [15:0] out_e3016;
wire  [15:0] out_e3017;
wire  [15:0] out_e3018;
wire  [15:0] out_e3019;
wire  [15:0] out_e3020;
wire  [15:0] out_e3021;
wire  [15:0] out_e3022;
wire  [15:0] out_e3023;
wire  [15:0] out_e3024;
wire  [15:0] out_e3025;
wire  [15:0] out_e3026;
wire  [15:0] out_e3027;
wire  [15:0] out_e3028;
wire  [15:0] out_e3029;
wire  [15:0] out_e3030;
wire  [15:0] out_e3031;
wire  [15:0] out_e3032;
wire  [15:0] out_e3033;
wire  [15:0] out_e3034;
wire  [15:0] out_e3035;
wire  [15:0] out_e3036;
wire  [15:0] out_e3037;
wire  [15:0] out_e3038;
wire  [15:0] out_e3039;
wire  [15:0] out_e3040;
wire  [15:0] out_e3041;
wire  [15:0] out_e3042;
wire  [15:0] out_e3043;
wire  [15:0] out_e3044;
wire  [15:0] out_e3045;
wire  [15:0] out_e3046;
wire  [15:0] out_e3047;
wire  [15:0] out_e3048;
wire  [15:0] out_e3049;
wire  [15:0] out_e3050;
wire  [15:0] out_e3051;
wire  [15:0] out_e3052;
wire  [15:0] out_e3053;
wire  [15:0] out_e3054;
wire  [15:0] out_e3055;
wire  [15:0] out_e3056;
wire  [15:0] out_e3057;
wire  [15:0] out_e3058;
wire  [15:0] out_e3059;
wire  [15:0] out_e3060;
wire  [15:0] out_e3061;
wire  [15:0] out_e3062;
wire  [15:0] out_e3063;
wire  [15:0] out_e3064;
wire  [15:0] out_e3065;
wire  [15:0] out_e3066;
wire  [15:0] out_e3067;
wire  [15:0] out_e3068;
wire  [15:0] out_e3069;
wire  [15:0] out_e3070;
wire  [15:0] out_e3071;
wire  [15:0] out_e3072;
wire  [15:0] out_e3073;
wire  [15:0] out_e3074;
wire  [15:0] out_e3075;
wire  [15:0] out_e3076;
wire  [15:0] out_e3077;
wire  [15:0] out_e3078;
wire  [15:0] out_e3079;
wire  [15:0] out_e3080;
wire  [15:0] out_e3081;
wire  [15:0] out_e3082;
wire  [15:0] out_e3083;
wire  [15:0] out_e3084;
wire  [15:0] out_e3085;
wire  [15:0] out_e3086;
wire  [15:0] out_e3087;
wire  [15:0] out_e3088;
wire  [15:0] out_e3089;
wire  [15:0] out_e3090;
wire  [15:0] out_e3091;
wire  [15:0] out_e3092;
wire  [15:0] out_e3093;
wire  [15:0] out_e3094;
wire  [15:0] out_e3095;
wire  [15:0] out_e3096;
wire  [15:0] out_e3097;
wire  [15:0] out_e3098;
wire  [15:0] out_e3099;
wire  [15:0] out_e3100;
wire  [15:0] out_e3101;
wire  [15:0] out_e3102;
wire  [15:0] out_e3103;
wire  [15:0] out_e3104;
wire  [15:0] out_e3105;
wire  [15:0] out_e3106;
wire  [15:0] out_e3107;
wire  [15:0] out_e3108;
wire  [15:0] out_e3109;
wire  [15:0] out_e3110;
wire  [15:0] out_e3111;
wire  [15:0] out_e3112;
wire  [15:0] out_e3113;
wire  [15:0] out_e3114;
wire  [15:0] out_e3115;
wire  [15:0] out_e3116;
wire  [15:0] out_e3117;
wire  [15:0] out_e3118;
wire  [15:0] out_e3119;
wire  [15:0] out_e3120;
wire  [15:0] out_e3121;
wire  [15:0] out_e3122;
wire  [15:0] out_e3123;
wire  [15:0] out_e3124;
wire  [15:0] out_e3125;
wire  [15:0] out_e3126;
wire  [15:0] out_e3127;
wire  [15:0] out_e3128;
wire  [15:0] out_e3129;
wire  [15:0] out_e3130;
wire  [15:0] out_e3131;
wire  [15:0] out_e3132;
wire  [15:0] out_e3133;
wire  [15:0] out_e3134;
wire  [15:0] out_e3135;
wire  [15:0] out_e3136;
wire  [15:0] out_e3137;
wire  [15:0] out_e3138;
wire  [15:0] out_e3139;
wire  [15:0] out_e3140;
wire  [15:0] out_e3141;
wire  [15:0] out_e3142;
wire  [15:0] out_e3143;
wire  [15:0] out_e3144;
wire  [15:0] out_e3145;
wire  [15:0] out_e3146;
wire  [15:0] out_e3147;
wire  [15:0] out_e3148;
wire  [15:0] out_e3149;
wire  [15:0] out_e3150;
wire  [15:0] out_e3151;
wire  [15:0] out_e3152;
wire  [15:0] out_e3153;
wire  [15:0] out_e3154;
wire  [15:0] out_e3155;
wire  [15:0] out_e3156;
wire  [15:0] out_e3157;
wire  [15:0] out_e3158;
wire  [15:0] out_e3159;
wire  [15:0] out_e3160;
wire  [15:0] out_e3161;
wire  [15:0] out_e3162;
wire  [15:0] out_e3163;
wire  [15:0] out_e3164;
wire  [15:0] out_e3165;
wire  [15:0] out_e3166;
wire  [15:0] out_e3167;
wire  [15:0] out_e3168;
wire  [15:0] out_e3169;
wire  [15:0] out_e3170;
wire  [15:0] out_e3171;
wire  [15:0] out_e3172;
wire  [15:0] out_e3173;
wire  [15:0] out_e3174;
wire  [15:0] out_e3175;
wire  [15:0] out_e3176;
wire  [15:0] out_e3177;
wire  [15:0] out_e3178;
wire  [15:0] out_e3179;
wire  [15:0] out_e3180;
wire  [15:0] out_e3181;
wire  [15:0] out_e3182;
wire  [15:0] out_e3183;
wire  [15:0] out_e3184;
wire  [15:0] out_e3185;
wire  [15:0] out_e3186;
wire  [15:0] out_e3187;
wire  [15:0] out_e3188;
wire  [15:0] out_e3189;
wire  [15:0] out_e3190;
wire  [15:0] out_e3191;
wire  [15:0] out_e3192;
wire  [15:0] out_e3193;
wire  [15:0] out_e3194;
wire  [15:0] out_e3195;
wire  [15:0] out_e3196;
wire  [15:0] out_e3197;
wire  [15:0] out_e3198;
wire  [15:0] out_e3199;
wire  [15:0] out_e3200;
wire  [15:0] out_e3201;
wire  [15:0] out_e3202;
wire  [15:0] out_e3203;
wire  [15:0] out_e3204;
wire  [15:0] out_e3205;
wire  [15:0] out_e3206;
wire  [15:0] out_e3207;
wire  [15:0] out_e3208;
wire  [15:0] out_e3209;
wire  [15:0] out_e3210;
wire  [15:0] out_e3211;
wire  [15:0] out_e3212;
wire  [15:0] out_e3213;
wire  [15:0] out_e3214;
wire  [15:0] out_e3215;
wire  [15:0] out_e3216;
wire  [15:0] out_e3217;
wire  [15:0] out_e3218;
wire  [15:0] out_e3219;
wire  [15:0] out_e3220;
wire  [15:0] out_e3221;
wire  [15:0] out_e3222;
wire  [15:0] out_e3223;
wire  [15:0] out_e3224;
wire  [15:0] out_e3225;
wire  [15:0] out_e3226;
wire  [15:0] out_e3227;
wire  [15:0] out_e3228;
wire  [15:0] out_e3229;
wire  [15:0] out_e3230;
wire  [15:0] out_e3231;
wire  [15:0] out_e3232;
wire  [15:0] out_e3233;
wire  [15:0] out_e3234;
wire  [15:0] out_e3235;
wire  [15:0] out_e3236;
wire  [15:0] out_e3237;
wire  [15:0] out_e3238;
wire  [15:0] out_e3239;
wire  [15:0] out_e3240;
wire  [15:0] out_e3241;
wire  [15:0] out_e3242;
wire  [15:0] out_e3243;
wire  [15:0] out_e3244;
wire  [15:0] out_e3245;
wire  [15:0] out_e3246;
wire  [15:0] out_e3247;
wire  [15:0] out_e3248;
wire  [15:0] out_e3249;
wire  [15:0] out_e3250;
wire  [15:0] out_e3251;
wire  [15:0] out_e3252;
wire  [15:0] out_e3253;
wire  [15:0] out_e3254;
wire  [15:0] out_e3255;
wire  [15:0] out_e3256;
wire  [15:0] out_e3257;
wire  [15:0] out_e3258;
wire  [15:0] out_e3259;
wire  [15:0] out_e3260;
wire  [15:0] out_e3261;
wire  [15:0] out_e3262;
wire  [15:0] out_e3263;
wire  [15:0] out_e3264;
wire  [15:0] out_e3265;
wire  [15:0] out_e3266;
wire  [15:0] out_e3267;
wire  [15:0] out_e3268;
wire  [15:0] out_e3269;
wire  [15:0] out_e3270;
wire  [15:0] out_e3271;
wire  [15:0] out_e3272;
wire  [15:0] out_e3273;
wire  [15:0] out_e3274;
wire  [15:0] out_e3275;
wire  [15:0] out_e3276;
wire  [15:0] out_e3277;
wire  [15:0] out_e3278;
wire  [15:0] out_e3279;
wire  [15:0] out_e3280;
wire  [15:0] out_e3281;
wire  [15:0] out_e3282;
wire  [15:0] out_e3283;
wire  [15:0] out_e3284;
wire  [15:0] out_e3285;
wire  [15:0] out_e3286;
wire  [15:0] out_e3287;
wire  [15:0] out_e3288;
wire  [15:0] out_e3289;
wire  [15:0] out_e3290;
wire  [15:0] out_e3291;
wire  [15:0] out_e3292;
wire  [15:0] out_e3293;
wire  [15:0] out_e3294;
wire  [15:0] out_e3295;
wire  [15:0] out_e3296;
wire  [15:0] out_e3297;
wire  [15:0] out_e3298;
wire  [15:0] out_e3299;
wire  [15:0] out_e3300;
wire  [15:0] out_e3301;
wire  [15:0] out_e3302;
wire  [15:0] out_e3303;
wire  [15:0] out_e3304;
wire  [15:0] out_e3305;
wire  [15:0] out_e3306;
wire  [15:0] out_e3307;
wire  [15:0] out_e3308;
wire  [15:0] out_e3309;
wire  [15:0] out_e3310;
wire  [15:0] out_e3311;
wire  [15:0] out_e3312;
wire  [15:0] out_e3313;
wire  [15:0] out_e3314;
wire  [15:0] out_e3315;
wire  [15:0] out_e3316;
wire  [15:0] out_e3317;
wire  [15:0] out_e3318;
wire  [15:0] out_e3319;
wire  [15:0] out_e3320;
wire  [15:0] out_e3321;
wire  [15:0] out_e3322;
wire  [15:0] out_e3323;
wire  [15:0] out_e3324;
wire  [15:0] out_e3325;
wire  [15:0] out_e3326;
wire  [15:0] out_e3327;
wire  [15:0] out_e3328;
wire  [15:0] out_e3329;
wire  [15:0] out_e3330;
wire  [15:0] out_e3331;
wire  [15:0] out_e3332;
wire  [15:0] out_e3333;
wire  [15:0] out_e3334;
wire  [15:0] out_e3335;
wire  [15:0] out_e3336;
wire  [15:0] out_e3337;
wire  [15:0] out_e3338;
wire  [15:0] out_e3339;
wire  [15:0] out_e3340;
wire  [15:0] out_e3341;
wire  [15:0] out_e3342;
wire  [15:0] out_e3343;
wire  [15:0] out_e3344;
wire  [15:0] out_e3345;
wire  [15:0] out_e3346;
wire  [15:0] out_e3347;
wire  [15:0] out_e3348;
wire  [15:0] out_e3349;
wire  [15:0] out_e3350;
wire  [15:0] out_e3351;
wire  [15:0] out_e3352;
wire  [15:0] out_e3353;
wire  [15:0] out_e3354;
wire  [15:0] out_e3355;
wire  [15:0] out_e3356;
wire  [15:0] out_e3357;
wire  [15:0] out_e3358;
wire  [15:0] out_e3359;
wire  [15:0] out_e3360;
wire  [15:0] out_e3361;
wire  [15:0] out_e3362;
wire  [15:0] out_e3363;
wire  [15:0] out_e3364;
wire  [15:0] out_e3365;
wire  [15:0] out_e3366;
wire  [15:0] out_e3367;
wire  [15:0] out_e3368;
wire  [15:0] out_e3369;
wire  [15:0] out_e3370;
wire  [15:0] out_e3371;
wire  [15:0] out_e3372;
wire  [15:0] out_e3373;
wire  [15:0] out_e3374;
wire  [15:0] out_e3375;
wire  [15:0] out_e3376;
wire  [15:0] out_e3377;
wire  [15:0] out_e3378;
wire  [15:0] out_e3379;
wire  [15:0] out_e3380;
wire  [15:0] out_e3381;
wire  [15:0] out_e3382;
wire  [15:0] out_e3383;
wire  [15:0] out_e3384;
wire  [15:0] out_e3385;
wire  [15:0] out_e3386;
wire  [15:0] out_e3387;
wire  [15:0] out_e3388;
wire  [15:0] out_e3389;
wire  [15:0] out_e3390;
wire  [15:0] out_e3391;
wire  [15:0] out_e3392;
wire  [15:0] out_e3393;
wire  [15:0] out_e3394;
wire  [15:0] out_e3395;
wire  [15:0] out_e3396;
wire  [15:0] out_e3397;
wire  [15:0] out_e3398;
wire  [15:0] out_e3399;
wire  [15:0] out_e3400;
wire  [15:0] out_e3401;
wire  [15:0] out_e3402;
wire  [15:0] out_e3403;
wire  [15:0] out_e3404;
wire  [15:0] out_e3405;
wire  [15:0] out_e3406;
wire  [15:0] out_e3407;
wire  [15:0] out_e3408;
wire  [15:0] out_e3409;
wire  [15:0] out_e3410;
wire  [15:0] out_e3411;
wire  [15:0] out_e3412;
wire  [15:0] out_e3413;
wire  [15:0] out_e3414;
wire  [15:0] out_e3415;
wire  [15:0] out_e3416;
wire  [15:0] out_e3417;
wire  [15:0] out_e3418;
wire  [15:0] out_e3419;
wire  [15:0] out_e3420;
wire  [15:0] out_e3421;
wire  [15:0] out_e3422;
wire  [15:0] out_e3423;
wire  [15:0] out_e3424;
wire  [15:0] out_e3425;
wire  [15:0] out_e3426;
wire  [15:0] out_e3427;
wire  [15:0] out_e3428;
wire  [15:0] out_e3429;
wire  [15:0] out_e3430;
wire  [15:0] out_e3431;
wire  [15:0] out_e3432;
wire  [15:0] out_e3433;
wire  [15:0] out_e3434;
wire  [15:0] out_e3435;
wire  [15:0] out_e3436;
wire  [15:0] out_e3437;
wire  [15:0] out_e3438;
wire  [15:0] out_e3439;
wire  [15:0] out_e3440;
wire  [15:0] out_e3441;
wire  [15:0] out_e3442;
wire  [15:0] out_e3443;
wire  [15:0] out_e3444;
wire  [15:0] out_e3445;
wire  [15:0] out_e3446;
wire  [15:0] out_e3447;
wire  [15:0] out_e3448;
wire  [15:0] out_e3449;
wire  [15:0] out_e3450;
wire  [15:0] out_e3451;
wire  [15:0] out_e3452;
wire  [15:0] out_e3453;
wire  [15:0] out_e3454;
wire  [15:0] out_e3455;
wire  [15:0] out_e3456;
wire  [15:0] out_e3457;
wire  [15:0] out_e3458;
wire  [15:0] out_e3459;
wire  [15:0] out_e3460;
wire  [15:0] out_e3461;
wire  [15:0] out_e3462;
wire  [15:0] out_e3463;
wire  [15:0] out_e3464;
wire  [15:0] out_e3465;
wire  [15:0] out_e3466;
wire  [15:0] out_e3467;
wire  [15:0] out_e3468;
wire  [15:0] out_e3469;
wire  [15:0] out_e3470;
wire  [15:0] out_e3471;
wire  [15:0] out_e3472;
wire  [15:0] out_e3473;
wire  [15:0] out_e3474;
wire  [15:0] out_e3475;
wire  [15:0] out_e3476;
wire  [15:0] out_e3477;
wire  [15:0] out_e3478;
wire  [15:0] out_e3479;
wire  [15:0] out_e3480;
wire  [15:0] out_e3481;
wire  [15:0] out_e3482;
wire  [15:0] out_e3483;
wire  [15:0] out_e3484;
wire  [15:0] out_e3485;
wire  [15:0] out_e3486;
wire  [15:0] out_e3487;
wire  [15:0] out_e3488;
wire  [15:0] out_e3489;
wire  [15:0] out_e3490;
wire  [15:0] out_e3491;
wire  [15:0] out_e3492;
wire  [15:0] out_e3493;
wire  [15:0] out_e3494;
wire  [15:0] out_e3495;
wire  [15:0] out_e3496;
wire  [15:0] out_e3497;
wire  [15:0] out_e3498;
wire  [15:0] out_e3499;
wire  [15:0] out_e3500;
wire  [15:0] out_e3501;
wire  [15:0] out_e3502;
wire  [15:0] out_e3503;
wire  [15:0] out_e3504;
wire  [15:0] out_e3505;
wire  [15:0] out_e3506;
wire  [15:0] out_e3507;
wire  [15:0] out_e3508;
wire  [15:0] out_e3509;
wire  [15:0] out_e3510;
wire  [15:0] out_e3511;
wire  [15:0] out_e3512;
wire  [15:0] out_e3513;
wire  [15:0] out_e3514;
wire  [15:0] out_e3515;
wire  [15:0] out_e3516;
wire  [15:0] out_e3517;
wire  [15:0] out_e3518;
wire  [15:0] out_e3519;
wire  [15:0] out_e3520;
wire  [15:0] out_e3521;
wire  [15:0] out_e3522;
wire  [15:0] out_e3523;
wire  [15:0] out_e3524;
wire  [15:0] out_e3525;
wire  [15:0] out_e3526;
wire  [15:0] out_e3527;
wire  [15:0] out_e3528;
wire  [15:0] out_e3529;
wire  [15:0] out_e3530;
wire  [15:0] out_e3531;
wire  [15:0] out_e3532;
wire  [15:0] out_e3533;
wire  [15:0] out_e3534;
wire  [15:0] out_e3535;
wire  [15:0] out_e3536;
wire  [15:0] out_e3537;
wire  [15:0] out_e3538;
wire  [15:0] out_e3539;
wire  [15:0] out_e3540;
wire  [15:0] out_e3541;
wire  [15:0] out_e3542;
wire  [15:0] out_e3543;
wire  [15:0] out_e3544;
wire  [15:0] out_e3545;
wire  [15:0] out_e3546;
wire  [15:0] out_e3547;
wire  [15:0] out_e3548;
wire  [15:0] out_e3549;
wire  [15:0] out_e3550;
wire  [15:0] out_e3551;
wire  [15:0] out_e3552;
wire  [15:0] out_e3553;
wire  [15:0] out_e3554;
wire  [15:0] out_e3555;
wire  [15:0] out_e3556;
wire  [15:0] out_e3557;
wire  [15:0] out_e3558;
wire  [15:0] out_e3559;
wire  [15:0] out_e3560;
wire  [15:0] out_e3561;
wire  [15:0] out_e3562;
wire  [15:0] out_e3563;
wire  [15:0] out_e3564;
wire  [15:0] out_e3565;
wire  [15:0] out_e3566;
wire  [15:0] out_e3567;
wire  [15:0] out_e3568;
wire  [15:0] out_e3569;
wire  [15:0] out_e3570;
wire  [15:0] out_e3571;
wire  [15:0] out_e3572;
wire  [15:0] out_e3573;
wire  [15:0] out_e3574;
wire  [15:0] out_e3575;
wire  [15:0] out_e3576;
wire  [15:0] out_e3577;
wire  [15:0] out_e3578;
wire  [15:0] out_e3579;
wire  [15:0] out_e3580;
wire  [15:0] out_e3581;
wire  [15:0] out_e3582;
wire  [15:0] out_e3583;
wire  [15:0] out_e3584;
wire  [15:0] out_e3585;
wire  [15:0] out_e3586;
wire  [15:0] out_e3587;
wire  [15:0] out_e3588;
wire  [15:0] out_e3589;
wire  [15:0] out_e3590;
wire  [15:0] out_e3591;
wire  [15:0] out_e3592;
wire  [15:0] out_e3593;
wire  [15:0] out_e3594;
wire  [15:0] out_e3595;
wire  [15:0] out_e3596;
wire  [15:0] out_e3597;
wire  [15:0] out_e3598;
wire  [15:0] out_e3599;
wire  [15:0] out_e3600;
wire  [15:0] out_e3601;
wire  [15:0] out_e3602;
wire  [15:0] out_e3603;
wire  [15:0] out_e3604;
wire  [15:0] out_e3605;
wire  [15:0] out_e3606;
wire  [15:0] out_e3607;
wire  [15:0] out_e3608;
wire  [15:0] out_e3609;
wire  [15:0] out_e3610;
wire  [15:0] out_e3611;
wire  [15:0] out_e3612;
wire  [15:0] out_e3613;
wire  [15:0] out_e3614;
wire  [15:0] out_e3615;
wire  [15:0] out_e3616;
wire  [15:0] out_e3617;
wire  [15:0] out_e3618;
wire  [15:0] out_e3619;
wire  [15:0] out_e3620;
wire  [15:0] out_e3621;
wire  [15:0] out_e3622;
wire  [15:0] out_e3623;
wire  [15:0] out_e3624;
wire  [15:0] out_e3625;
wire  [15:0] out_e3626;
wire  [15:0] out_e3627;
wire  [15:0] out_e3628;
wire  [15:0] out_e3629;
wire  [15:0] out_e3630;
wire  [15:0] out_e3631;
wire  [15:0] out_e3632;
wire  [15:0] out_e3633;
wire  [15:0] out_e3634;
wire  [15:0] out_e3635;
wire  [15:0] out_e3636;
wire  [15:0] out_e3637;
wire  [15:0] out_e3638;
wire  [15:0] out_e3639;
wire  [15:0] out_e3640;
wire  [15:0] out_e3641;
wire  [15:0] out_e3642;
wire  [15:0] out_e3643;
wire  [15:0] out_e3644;
wire  [15:0] out_e3645;
wire  [15:0] out_e3646;
wire  [15:0] out_e3647;
wire  [15:0] out_e3648;
wire  [15:0] out_e3649;
wire  [15:0] out_e3650;
wire  [15:0] out_e3651;
wire  [15:0] out_e3652;
wire  [15:0] out_e3653;
wire  [15:0] out_e3654;
wire  [15:0] out_e3655;
wire  [15:0] out_e3656;
wire  [15:0] out_e3657;
wire  [15:0] out_e3658;
wire  [15:0] out_e3659;
wire  [15:0] out_e3660;
wire  [15:0] out_e3661;
wire  [15:0] out_e3662;
wire  [15:0] out_e3663;
wire  [15:0] out_e3664;
wire  [15:0] out_e3665;
wire  [15:0] out_e3666;
wire  [15:0] out_e3667;
wire  [15:0] out_e3668;
wire  [15:0] out_e3669;
wire  [15:0] out_e3670;
wire  [15:0] out_e3671;
wire  [15:0] out_e3672;
wire  [15:0] out_e3673;
wire  [15:0] out_e3674;
wire  [15:0] out_e3675;
wire  [15:0] out_e3676;
wire  [15:0] out_e3677;
wire  [15:0] out_e3678;
wire  [15:0] out_e3679;
wire  [15:0] out_e3680;
wire  [15:0] out_e3681;
wire  [15:0] out_e3682;
wire  [15:0] out_e3683;
wire  [15:0] out_e3684;
wire  [15:0] out_e3685;
wire  [15:0] out_e3686;
wire  [15:0] out_e3687;
wire  [15:0] out_e3688;
wire  [15:0] out_e3689;
wire  [15:0] out_e3690;
wire  [15:0] out_e3691;
wire  [15:0] out_e3692;
wire  [15:0] out_e3693;
wire  [15:0] out_e3694;
wire  [15:0] out_e3695;
wire  [15:0] out_e3696;
wire  [15:0] out_e3697;
wire  [15:0] out_e3698;
wire  [15:0] out_e3699;
wire  [15:0] out_e3700;
wire  [15:0] out_e3701;
wire  [15:0] out_e3702;
wire  [15:0] out_e3703;
wire  [15:0] out_e3704;
wire  [15:0] out_e3705;
wire  [15:0] out_e3706;
wire  [15:0] out_e3707;
wire  [15:0] out_e3708;
wire  [15:0] out_e3709;
wire  [15:0] out_e3710;
wire  [15:0] out_e3711;
wire  [15:0] out_e3712;
wire  [15:0] out_e3713;
wire  [15:0] out_e3714;
wire  [15:0] out_e3715;
wire  [15:0] out_e3716;
wire  [15:0] out_e3717;
wire  [15:0] out_e3718;
wire  [15:0] out_e3719;
wire  [15:0] out_e3720;
wire  [15:0] out_e3721;
wire  [15:0] out_e3722;
wire  [15:0] out_e3723;
wire  [15:0] out_e3724;
wire  [15:0] out_e3725;
wire  [15:0] out_e3726;
wire  [15:0] out_e3727;
wire  [15:0] out_e3728;
wire  [15:0] out_e3729;
wire  [15:0] out_e3730;
wire  [15:0] out_e3731;
wire  [15:0] out_e3732;
wire  [15:0] out_e3733;
wire  [15:0] out_e3734;
wire  [15:0] out_e3735;
wire  [15:0] out_e3736;
wire  [15:0] out_e3737;
wire  [15:0] out_e3738;
wire  [15:0] out_e3739;
wire  [15:0] out_e3740;
wire  [15:0] out_e3741;
wire  [15:0] out_e3742;
wire  [15:0] out_e3743;
wire  [15:0] out_e3744;
wire  [15:0] out_e3745;
wire  [15:0] out_e3746;
wire  [15:0] out_e3747;
wire  [15:0] out_e3748;
wire  [15:0] out_e3749;
wire  [15:0] out_e3750;
wire  [15:0] out_e3751;
wire  [15:0] out_e3752;
wire  [15:0] out_e3753;
wire  [15:0] out_e3754;
wire  [15:0] out_e3755;
wire  [15:0] out_e3756;
wire  [15:0] out_e3757;
wire  [15:0] out_e3758;
wire  [15:0] out_e3759;
wire  [15:0] out_e3760;
wire  [15:0] out_e3761;
wire  [15:0] out_e3762;
wire  [15:0] out_e3763;
wire  [15:0] out_e3764;
wire  [15:0] out_e3765;
wire  [15:0] out_e3766;
wire  [15:0] out_e3767;
wire  [15:0] out_e3768;
wire  [15:0] out_e3769;
wire  [15:0] out_e3770;
wire  [15:0] out_e3771;
wire  [15:0] out_e3772;
wire  [15:0] out_e3773;
wire  [15:0] out_e3774;
wire  [15:0] out_e3775;
wire  [15:0] out_e3776;
wire  [15:0] out_e3777;
wire  [15:0] out_e3778;
wire  [15:0] out_e3779;
wire  [15:0] out_e3780;
wire  [15:0] out_e3781;
wire  [15:0] out_e3782;
wire  [15:0] out_e3783;
wire  [15:0] out_e3784;
wire  [15:0] out_e3785;
wire  [15:0] out_e3786;
wire  [15:0] out_e3787;
wire  [15:0] out_e3788;
wire  [15:0] out_e3789;
wire  [15:0] out_e3790;
wire  [15:0] out_e3791;
wire  [15:0] out_e3792;
wire  [15:0] out_e3793;
wire  [15:0] out_e3794;
wire  [15:0] out_e3795;
wire  [15:0] out_e3796;
wire  [15:0] out_e3797;
wire  [15:0] out_e3798;
wire  [15:0] out_e3799;
wire  [15:0] out_e3800;
wire  [15:0] out_e3801;
wire  [15:0] out_e3802;
wire  [15:0] out_e3803;
wire  [15:0] out_e3804;
wire  [15:0] out_e3805;
wire  [15:0] out_e3806;
wire  [15:0] out_e3807;
wire  [15:0] out_e3808;
wire  [15:0] out_e3809;
wire  [15:0] out_e3810;
wire  [15:0] out_e3811;
wire  [15:0] out_e3812;
wire  [15:0] out_e3813;
wire  [15:0] out_e3814;
wire  [15:0] out_e3815;
wire  [15:0] out_e3816;
wire  [15:0] out_e3817;
wire  [15:0] out_e3818;
wire  [15:0] out_e3819;
wire  [15:0] out_e3820;
wire  [15:0] out_e3821;
wire  [15:0] out_e3822;
wire  [15:0] out_e3823;
wire  [15:0] out_e3824;
wire  [15:0] out_e3825;
wire  [15:0] out_e3826;
wire  [15:0] out_e3827;
wire  [15:0] out_e3828;
wire  [15:0] out_e3829;
wire  [15:0] out_e3830;
wire  [15:0] out_e3831;
wire  [15:0] out_e3832;
wire  [15:0] out_e3833;
wire  [15:0] out_e3834;
wire  [15:0] out_e3835;
wire  [15:0] out_e3836;
wire  [15:0] out_e3837;
wire  [15:0] out_e3838;
wire  [15:0] out_e3839;
wire  [15:0] out_e3840;
wire  [15:0] out_e3841;
wire  [15:0] out_e3842;
wire  [15:0] out_e3843;
wire  [15:0] out_e3844;
wire  [15:0] out_e3845;
wire  [15:0] out_e3846;
wire  [15:0] out_e3847;
wire  [15:0] out_e3848;
wire  [15:0] out_e3849;
wire  [15:0] out_e3850;
wire  [15:0] out_e3851;
wire  [15:0] out_e3852;
wire  [15:0] out_e3853;
wire  [15:0] out_e3854;
wire  [15:0] out_e3855;
wire  [15:0] out_e3856;
wire  [15:0] out_e3857;
wire  [15:0] out_e3858;
wire  [15:0] out_e3859;
wire  [15:0] out_e3860;
wire  [15:0] out_e3861;
wire  [15:0] out_e3862;
wire  [15:0] out_e3863;
wire  [15:0] out_e3864;
wire  [15:0] out_e3865;
wire  [15:0] out_e3866;
wire  [15:0] out_e3867;
wire  [15:0] out_e3868;
wire  [15:0] out_e3869;
wire  [15:0] out_e3870;
wire  [15:0] out_e3871;
wire  [15:0] out_e3872;
wire  [15:0] out_e3873;
wire  [15:0] out_e3874;
wire  [15:0] out_e3875;
wire  [15:0] out_e3876;
wire  [15:0] out_e3877;
wire  [15:0] out_e3878;
wire  [15:0] out_e3879;
wire  [15:0] out_e3880;
wire  [15:0] out_e3881;
wire  [15:0] out_e3882;
wire  [15:0] out_e3883;
wire  [15:0] out_e3884;
wire  [15:0] out_e3885;
wire  [15:0] out_e3886;
wire  [15:0] out_e3887;
wire  [15:0] out_e3888;
wire  [15:0] out_e3889;
wire  [15:0] out_e3890;
wire  [15:0] out_e3891;
wire  [15:0] out_e3892;
wire  [15:0] out_e3893;
wire  [15:0] out_e3894;
wire  [15:0] out_e3895;
wire  [15:0] out_e3896;
wire  [15:0] out_e3897;
wire  [15:0] out_e3898;
wire  [15:0] out_e3899;
wire  [15:0] out_e3900;
wire  [15:0] out_e3901;
wire  [15:0] out_e3902;
wire  [15:0] out_e3903;
wire  [15:0] out_e3904;
wire  [15:0] out_e3905;
wire  [15:0] out_e3906;
wire  [15:0] out_e3907;
wire  [15:0] out_e3908;
wire  [15:0] out_e3909;
wire  [15:0] out_e3910;
wire  [15:0] out_e3911;
wire  [15:0] out_e3912;
wire  [15:0] out_e3913;
wire  [15:0] out_e3914;
wire  [15:0] out_e3915;
wire  [15:0] out_e3916;
wire  [15:0] out_e3917;
wire  [15:0] out_e3918;
wire  [15:0] out_e3919;
wire  [15:0] out_e3920;
wire  [15:0] out_e3921;
wire  [15:0] out_e3922;
wire  [15:0] out_e3923;
wire  [15:0] out_e3924;
wire  [15:0] out_e3925;
wire  [15:0] out_e3926;
wire  [15:0] out_e3927;
wire  [15:0] out_e3928;
wire  [15:0] out_e3929;
wire  [15:0] out_e3930;
wire  [15:0] out_e3931;
wire  [15:0] out_e3932;
wire  [15:0] out_e3933;
wire  [15:0] out_e3934;
wire  [15:0] out_e3935;
wire  [15:0] out_e3936;
wire  [15:0] out_e3937;
wire  [15:0] out_e3938;
wire  [15:0] out_e3939;
wire  [15:0] out_e3940;
wire  [15:0] out_e3941;
wire  [15:0] out_e3942;
wire  [15:0] out_e3943;
wire  [15:0] out_e3944;
wire  [15:0] out_e3945;
wire  [15:0] out_e3946;
wire  [15:0] out_e3947;
wire  [15:0] out_e3948;
wire  [15:0] out_e3949;
wire  [15:0] out_e3950;
wire  [15:0] out_e3951;
wire  [15:0] out_e3952;
wire  [15:0] out_e3953;
wire  [15:0] out_e3954;
wire  [15:0] out_e3955;
wire  [15:0] out_e3956;
wire  [15:0] out_e3957;
wire  [15:0] out_e3958;
wire  [15:0] out_e3959;
wire  [15:0] out_e3960;
wire  [15:0] out_e3961;
wire  [15:0] out_e3962;
wire  [15:0] out_e3963;
wire  [15:0] out_e3964;
wire  [15:0] out_e3965;
wire  [15:0] out_e3966;
wire  [15:0] out_e3967;
wire  [15:0] out_e3968;
wire  [15:0] out_e3969;
wire  [15:0] out_e3970;
wire  [15:0] out_e3971;
wire  [15:0] out_e3972;
wire  [15:0] out_e3973;
wire  [15:0] out_e3974;
wire  [15:0] out_e3975;
wire  [15:0] out_e3976;
wire  [15:0] out_e3977;
wire  [15:0] out_e3978;
wire  [15:0] out_e3979;
wire  [15:0] out_e3980;
wire  [15:0] out_e3981;
wire  [15:0] out_e3982;
wire  [15:0] out_e3983;
wire  [15:0] out_e3984;
wire  [15:0] out_e3985;
wire  [15:0] out_e3986;
wire  [15:0] out_e3987;
wire  [15:0] out_e3988;
wire  [15:0] out_e3989;
wire  [15:0] out_e3990;
wire  [15:0] out_e3991;
wire  [15:0] out_e3992;
wire  [15:0] out_e3993;
wire  [15:0] out_e3994;
wire  [15:0] out_e3995;
wire  [15:0] out_e3996;
wire  [15:0] out_e3997;
wire  [15:0] out_e3998;
wire  [15:0] out_e3999;
wire  [15:0] out_e4000;
wire  [15:0] out_e4001;
wire  [15:0] out_e4002;
wire  [15:0] out_e4003;
wire  [15:0] out_e4004;
wire  [15:0] out_e4005;
wire  [15:0] out_e4006;
wire  [15:0] out_e4007;
wire  [15:0] out_e4008;
wire  [15:0] out_e4009;
wire  [15:0] out_e4010;
wire  [15:0] out_e4011;
wire  [15:0] out_e4012;
wire  [15:0] out_e4013;
wire  [15:0] out_e4014;
wire  [15:0] out_e4015;
wire  [15:0] out_e4016;
wire  [15:0] out_e4017;
wire  [15:0] out_e4018;
wire  [15:0] out_e4019;
wire  [15:0] out_e4020;
wire  [15:0] out_e4021;
wire  [15:0] out_e4022;
wire  [15:0] out_e4023;
wire  [15:0] out_e4024;
wire  [15:0] out_e4025;
wire  [15:0] out_e4026;
wire  [15:0] out_e4027;
wire  [15:0] out_e4028;
wire  [15:0] out_e4029;
wire  [15:0] out_e4030;
wire  [15:0] out_e4031;
wire  [15:0] out_e4032;
wire  [15:0] out_e4033;
wire  [15:0] out_e4034;
wire  [15:0] out_e4035;
wire  [15:0] out_e4036;
wire  [15:0] out_e4037;
wire  [15:0] out_e4038;
wire  [15:0] out_e4039;
wire  [15:0] out_e4040;
wire  [15:0] out_e4041;
wire  [15:0] out_e4042;
wire  [15:0] out_e4043;
wire  [15:0] out_e4044;
wire  [15:0] out_e4045;
wire  [15:0] out_e4046;
wire  [15:0] out_e4047;
wire  [15:0] out_e4048;
wire  [15:0] out_e4049;
wire  [15:0] out_e4050;
wire  [15:0] out_e4051;
wire  [15:0] out_e4052;
wire  [15:0] out_e4053;
wire  [15:0] out_e4054;
wire  [15:0] out_e4055;
wire  [15:0] out_e4056;
wire  [15:0] out_e4057;
wire  [15:0] out_e4058;
wire  [15:0] out_e4059;
wire  [15:0] out_e4060;
wire  [15:0] out_e4061;
wire  [15:0] out_e4062;
wire  [15:0] out_e4063;
wire  [15:0] out_e4064;
wire  [15:0] out_e4065;
wire  [15:0] out_e4066;
wire  [15:0] out_e4067;
wire  [15:0] out_e4068;
wire  [15:0] out_e4069;
wire  [15:0] out_e4070;
wire  [15:0] out_e4071;
wire  [15:0] out_e4072;
wire  [15:0] out_e4073;
wire  [15:0] out_e4074;
wire  [15:0] out_e4075;
wire  [15:0] out_e4076;
wire  [15:0] out_e4077;
wire  [15:0] out_e4078;
wire  [15:0] out_e4079;
wire  [15:0] out_e4080;
wire  [15:0] out_e4081;
wire  [15:0] out_e4082;
wire  [15:0] out_e4083;
wire  [15:0] out_e4084;
wire  [15:0] out_e4085;
wire  [15:0] out_e4086;
wire  [15:0] out_e4087;
wire  [15:0] out_e4088;
wire  [15:0] out_e4089;
wire  [15:0] out_e4090;
wire  [15:0] out_e4091;
wire  [15:0] out_e4092;
wire  [15:0] out_e4093;
wire  [15:0] out_e4094;
wire  [15:0] out_e4095;

wire  [15:0] result0;
wire  [15:0] result1;
wire  [15:0] result2;
wire  [15:0] result3;
wire  [15:0] result4;
wire  [15:0] result5;
wire  [15:0] result6;
wire  [15:0] result7;
wire  [15:0] result8;
wire  [15:0] result9;
wire  [15:0] result10;
wire  [15:0] result11;
wire  [15:0] result12;
wire  [15:0] result13;
wire  [15:0] result14;
wire  [15:0] result15;
wire  [15:0] result16;
wire  [15:0] result17;
wire  [15:0] result18;
wire  [15:0] result19;
wire  [15:0] result20;
wire  [15:0] result21;
wire  [15:0] result22;
wire  [15:0] result23;
wire  [15:0] result24;
wire  [15:0] result25;
wire  [15:0] result26;
wire  [15:0] result27;
wire  [15:0] result28;
wire  [15:0] result29;
wire  [15:0] result30;
wire  [15:0] result31;
wire  [15:0] result32;
wire  [15:0] result33;
wire  [15:0] result34;
wire  [15:0] result35;
wire  [15:0] result36;
wire  [15:0] result37;
wire  [15:0] result38;
wire  [15:0] result39;
wire  [15:0] result40;
wire  [15:0] result41;
wire  [15:0] result42;
wire  [15:0] result43;
wire  [15:0] result44;
wire  [15:0] result45;
wire  [15:0] result46;
wire  [15:0] result47;
wire  [15:0] result48;
wire  [15:0] result49;
wire  [15:0] result50;
wire  [15:0] result51;
wire  [15:0] result52;
wire  [15:0] result53;
wire  [15:0] result54;
wire  [15:0] result55;
wire  [15:0] result56;
wire  [15:0] result57;
wire  [15:0] result58;
wire  [15:0] result59;
wire  [15:0] result60;
wire  [15:0] result61;
wire  [15:0] result62;
wire  [15:0] result63;
wire  [15:0] result64;
wire  [15:0] result65;
wire  [15:0] result66;
wire  [15:0] result67;
wire  [15:0] result68;
wire  [15:0] result69;
wire  [15:0] result70;
wire  [15:0] result71;
wire  [15:0] result72;
wire  [15:0] result73;
wire  [15:0] result74;
wire  [15:0] result75;
wire  [15:0] result76;
wire  [15:0] result77;
wire  [15:0] result78;
wire  [15:0] result79;
wire  [15:0] result80;
wire  [15:0] result81;
wire  [15:0] result82;
wire  [15:0] result83;
wire  [15:0] result84;
wire  [15:0] result85;
wire  [15:0] result86;
wire  [15:0] result87;
wire  [15:0] result88;
wire  [15:0] result89;
wire  [15:0] result90;
wire  [15:0] result91;
wire  [15:0] result92;
wire  [15:0] result93;
wire  [15:0] result94;
wire  [15:0] result95;
wire  [15:0] result96;
wire  [15:0] result97;
wire  [15:0] result98;
wire  [15:0] result99;
wire  [15:0] result100;
wire  [15:0] result101;
wire  [15:0] result102;
wire  [15:0] result103;
wire  [15:0] result104;
wire  [15:0] result105;
wire  [15:0] result106;
wire  [15:0] result107;
wire  [15:0] result108;
wire  [15:0] result109;
wire  [15:0] result110;
wire  [15:0] result111;
wire  [15:0] result112;
wire  [15:0] result113;
wire  [15:0] result114;
wire  [15:0] result115;
wire  [15:0] result116;
wire  [15:0] result117;
wire  [15:0] result118;
wire  [15:0] result119;
wire  [15:0] result120;
wire  [15:0] result121;
wire  [15:0] result122;
wire  [15:0] result123;
wire  [15:0] result124;
wire  [15:0] result125;
wire  [15:0] result126;
wire  [15:0] result127;
wire  [15:0] result128;
wire  [15:0] result129;
wire  [15:0] result130;
wire  [15:0] result131;
wire  [15:0] result132;
wire  [15:0] result133;
wire  [15:0] result134;
wire  [15:0] result135;
wire  [15:0] result136;
wire  [15:0] result137;
wire  [15:0] result138;
wire  [15:0] result139;
wire  [15:0] result140;
wire  [15:0] result141;
wire  [15:0] result142;
wire  [15:0] result143;
wire  [15:0] result144;
wire  [15:0] result145;
wire  [15:0] result146;
wire  [15:0] result147;
wire  [15:0] result148;
wire  [15:0] result149;
wire  [15:0] result150;
wire  [15:0] result151;
wire  [15:0] result152;
wire  [15:0] result153;
wire  [15:0] result154;
wire  [15:0] result155;
wire  [15:0] result156;
wire  [15:0] result157;
wire  [15:0] result158;
wire  [15:0] result159;
wire  [15:0] result160;
wire  [15:0] result161;
wire  [15:0] result162;
wire  [15:0] result163;
wire  [15:0] result164;
wire  [15:0] result165;
wire  [15:0] result166;
wire  [15:0] result167;
wire  [15:0] result168;
wire  [15:0] result169;
wire  [15:0] result170;
wire  [15:0] result171;
wire  [15:0] result172;
wire  [15:0] result173;
wire  [15:0] result174;
wire  [15:0] result175;
wire  [15:0] result176;
wire  [15:0] result177;
wire  [15:0] result178;
wire  [15:0] result179;
wire  [15:0] result180;
wire  [15:0] result181;
wire  [15:0] result182;
wire  [15:0] result183;
wire  [15:0] result184;
wire  [15:0] result185;
wire  [15:0] result186;
wire  [15:0] result187;
wire  [15:0] result188;
wire  [15:0] result189;
wire  [15:0] result190;
wire  [15:0] result191;
wire  [15:0] result192;
wire  [15:0] result193;
wire  [15:0] result194;
wire  [15:0] result195;
wire  [15:0] result196;
wire  [15:0] result197;
wire  [15:0] result198;
wire  [15:0] result199;
wire  [15:0] result200;
wire  [15:0] result201;
wire  [15:0] result202;
wire  [15:0] result203;
wire  [15:0] result204;
wire  [15:0] result205;
wire  [15:0] result206;
wire  [15:0] result207;
wire  [15:0] result208;
wire  [15:0] result209;
wire  [15:0] result210;
wire  [15:0] result211;
wire  [15:0] result212;
wire  [15:0] result213;
wire  [15:0] result214;
wire  [15:0] result215;
wire  [15:0] result216;
wire  [15:0] result217;
wire  [15:0] result218;
wire  [15:0] result219;
wire  [15:0] result220;
wire  [15:0] result221;
wire  [15:0] result222;
wire  [15:0] result223;
wire  [15:0] result224;
wire  [15:0] result225;
wire  [15:0] result226;
wire  [15:0] result227;
wire  [15:0] result228;
wire  [15:0] result229;
wire  [15:0] result230;
wire  [15:0] result231;
wire  [15:0] result232;
wire  [15:0] result233;
wire  [15:0] result234;
wire  [15:0] result235;
wire  [15:0] result236;
wire  [15:0] result237;
wire  [15:0] result238;
wire  [15:0] result239;
wire  [15:0] result240;
wire  [15:0] result241;
wire  [15:0] result242;
wire  [15:0] result243;
wire  [15:0] result244;
wire  [15:0] result245;
wire  [15:0] result246;
wire  [15:0] result247;
wire  [15:0] result248;
wire  [15:0] result249;
wire  [15:0] result250;
wire  [15:0] result251;
wire  [15:0] result252;
wire  [15:0] result253;
wire  [15:0] result254;
wire  [15:0] result255;
wire  [15:0] result256;
wire  [15:0] result257;
wire  [15:0] result258;
wire  [15:0] result259;
wire  [15:0] result260;
wire  [15:0] result261;
wire  [15:0] result262;
wire  [15:0] result263;
wire  [15:0] result264;
wire  [15:0] result265;
wire  [15:0] result266;
wire  [15:0] result267;
wire  [15:0] result268;
wire  [15:0] result269;
wire  [15:0] result270;
wire  [15:0] result271;
wire  [15:0] result272;
wire  [15:0] result273;
wire  [15:0] result274;
wire  [15:0] result275;
wire  [15:0] result276;
wire  [15:0] result277;
wire  [15:0] result278;
wire  [15:0] result279;
wire  [15:0] result280;
wire  [15:0] result281;
wire  [15:0] result282;
wire  [15:0] result283;
wire  [15:0] result284;
wire  [15:0] result285;
wire  [15:0] result286;
wire  [15:0] result287;
wire  [15:0] result288;
wire  [15:0] result289;
wire  [15:0] result290;
wire  [15:0] result291;
wire  [15:0] result292;
wire  [15:0] result293;
wire  [15:0] result294;
wire  [15:0] result295;
wire  [15:0] result296;
wire  [15:0] result297;
wire  [15:0] result298;
wire  [15:0] result299;
wire  [15:0] result300;
wire  [15:0] result301;
wire  [15:0] result302;
wire  [15:0] result303;
wire  [15:0] result304;
wire  [15:0] result305;
wire  [15:0] result306;
wire  [15:0] result307;
wire  [15:0] result308;
wire  [15:0] result309;
wire  [15:0] result310;
wire  [15:0] result311;
wire  [15:0] result312;
wire  [15:0] result313;
wire  [15:0] result314;
wire  [15:0] result315;
wire  [15:0] result316;
wire  [15:0] result317;
wire  [15:0] result318;
wire  [15:0] result319;
wire  [15:0] result320;
wire  [15:0] result321;
wire  [15:0] result322;
wire  [15:0] result323;
wire  [15:0] result324;
wire  [15:0] result325;
wire  [15:0] result326;
wire  [15:0] result327;
wire  [15:0] result328;
wire  [15:0] result329;
wire  [15:0] result330;
wire  [15:0] result331;
wire  [15:0] result332;
wire  [15:0] result333;
wire  [15:0] result334;
wire  [15:0] result335;
wire  [15:0] result336;
wire  [15:0] result337;
wire  [15:0] result338;
wire  [15:0] result339;
wire  [15:0] result340;
wire  [15:0] result341;
wire  [15:0] result342;
wire  [15:0] result343;
wire  [15:0] result344;
wire  [15:0] result345;
wire  [15:0] result346;
wire  [15:0] result347;
wire  [15:0] result348;
wire  [15:0] result349;
wire  [15:0] result350;
wire  [15:0] result351;
wire  [15:0] result352;
wire  [15:0] result353;
wire  [15:0] result354;
wire  [15:0] result355;
wire  [15:0] result356;
wire  [15:0] result357;
wire  [15:0] result358;
wire  [15:0] result359;
wire  [15:0] result360;
wire  [15:0] result361;
wire  [15:0] result362;
wire  [15:0] result363;
wire  [15:0] result364;
wire  [15:0] result365;
wire  [15:0] result366;
wire  [15:0] result367;
wire  [15:0] result368;
wire  [15:0] result369;
wire  [15:0] result370;
wire  [15:0] result371;
wire  [15:0] result372;
wire  [15:0] result373;
wire  [15:0] result374;
wire  [15:0] result375;
wire  [15:0] result376;
wire  [15:0] result377;
wire  [15:0] result378;
wire  [15:0] result379;
wire  [15:0] result380;
wire  [15:0] result381;
wire  [15:0] result382;
wire  [15:0] result383;
wire  [15:0] result384;
wire  [15:0] result385;
wire  [15:0] result386;
wire  [15:0] result387;
wire  [15:0] result388;
wire  [15:0] result389;
wire  [15:0] result390;
wire  [15:0] result391;
wire  [15:0] result392;
wire  [15:0] result393;
wire  [15:0] result394;
wire  [15:0] result395;
wire  [15:0] result396;
wire  [15:0] result397;
wire  [15:0] result398;
wire  [15:0] result399;
wire  [15:0] result400;
wire  [15:0] result401;
wire  [15:0] result402;
wire  [15:0] result403;
wire  [15:0] result404;
wire  [15:0] result405;
wire  [15:0] result406;
wire  [15:0] result407;
wire  [15:0] result408;
wire  [15:0] result409;
wire  [15:0] result410;
wire  [15:0] result411;
wire  [15:0] result412;
wire  [15:0] result413;
wire  [15:0] result414;
wire  [15:0] result415;
wire  [15:0] result416;
wire  [15:0] result417;
wire  [15:0] result418;
wire  [15:0] result419;
wire  [15:0] result420;
wire  [15:0] result421;
wire  [15:0] result422;
wire  [15:0] result423;
wire  [15:0] result424;
wire  [15:0] result425;
wire  [15:0] result426;
wire  [15:0] result427;
wire  [15:0] result428;
wire  [15:0] result429;
wire  [15:0] result430;
wire  [15:0] result431;
wire  [15:0] result432;
wire  [15:0] result433;
wire  [15:0] result434;
wire  [15:0] result435;
wire  [15:0] result436;
wire  [15:0] result437;
wire  [15:0] result438;
wire  [15:0] result439;
wire  [15:0] result440;
wire  [15:0] result441;
wire  [15:0] result442;
wire  [15:0] result443;
wire  [15:0] result444;
wire  [15:0] result445;
wire  [15:0] result446;
wire  [15:0] result447;
wire  [15:0] result448;
wire  [15:0] result449;
wire  [15:0] result450;
wire  [15:0] result451;
wire  [15:0] result452;
wire  [15:0] result453;
wire  [15:0] result454;
wire  [15:0] result455;
wire  [15:0] result456;
wire  [15:0] result457;
wire  [15:0] result458;
wire  [15:0] result459;
wire  [15:0] result460;
wire  [15:0] result461;
wire  [15:0] result462;
wire  [15:0] result463;
wire  [15:0] result464;
wire  [15:0] result465;
wire  [15:0] result466;
wire  [15:0] result467;
wire  [15:0] result468;
wire  [15:0] result469;
wire  [15:0] result470;
wire  [15:0] result471;
wire  [15:0] result472;
wire  [15:0] result473;
wire  [15:0] result474;
wire  [15:0] result475;
wire  [15:0] result476;
wire  [15:0] result477;
wire  [15:0] result478;
wire  [15:0] result479;
wire  [15:0] result480;
wire  [15:0] result481;
wire  [15:0] result482;
wire  [15:0] result483;
wire  [15:0] result484;
wire  [15:0] result485;
wire  [15:0] result486;
wire  [15:0] result487;
wire  [15:0] result488;
wire  [15:0] result489;
wire  [15:0] result490;
wire  [15:0] result491;
wire  [15:0] result492;
wire  [15:0] result493;
wire  [15:0] result494;
wire  [15:0] result495;
wire  [15:0] result496;
wire  [15:0] result497;
wire  [15:0] result498;
wire  [15:0] result499;
wire  [15:0] result500;
wire  [15:0] result501;
wire  [15:0] result502;
wire  [15:0] result503;
wire  [15:0] result504;
wire  [15:0] result505;
wire  [15:0] result506;
wire  [15:0] result507;
wire  [15:0] result508;
wire  [15:0] result509;
wire  [15:0] result510;
wire  [15:0] result511;
wire  [15:0] result512;
wire  [15:0] result513;
wire  [15:0] result514;
wire  [15:0] result515;
wire  [15:0] result516;
wire  [15:0] result517;
wire  [15:0] result518;
wire  [15:0] result519;
wire  [15:0] result520;
wire  [15:0] result521;
wire  [15:0] result522;
wire  [15:0] result523;
wire  [15:0] result524;
wire  [15:0] result525;
wire  [15:0] result526;
wire  [15:0] result527;
wire  [15:0] result528;
wire  [15:0] result529;
wire  [15:0] result530;
wire  [15:0] result531;
wire  [15:0] result532;
wire  [15:0] result533;
wire  [15:0] result534;
wire  [15:0] result535;
wire  [15:0] result536;
wire  [15:0] result537;
wire  [15:0] result538;
wire  [15:0] result539;
wire  [15:0] result540;
wire  [15:0] result541;
wire  [15:0] result542;
wire  [15:0] result543;
wire  [15:0] result544;
wire  [15:0] result545;
wire  [15:0] result546;
wire  [15:0] result547;
wire  [15:0] result548;
wire  [15:0] result549;
wire  [15:0] result550;
wire  [15:0] result551;
wire  [15:0] result552;
wire  [15:0] result553;
wire  [15:0] result554;
wire  [15:0] result555;
wire  [15:0] result556;
wire  [15:0] result557;
wire  [15:0] result558;
wire  [15:0] result559;
wire  [15:0] result560;
wire  [15:0] result561;
wire  [15:0] result562;
wire  [15:0] result563;
wire  [15:0] result564;
wire  [15:0] result565;
wire  [15:0] result566;
wire  [15:0] result567;
wire  [15:0] result568;
wire  [15:0] result569;
wire  [15:0] result570;
wire  [15:0] result571;
wire  [15:0] result572;
wire  [15:0] result573;
wire  [15:0] result574;
wire  [15:0] result575;
wire  [15:0] result576;
wire  [15:0] result577;
wire  [15:0] result578;
wire  [15:0] result579;
wire  [15:0] result580;
wire  [15:0] result581;
wire  [15:0] result582;
wire  [15:0] result583;
wire  [15:0] result584;
wire  [15:0] result585;
wire  [15:0] result586;
wire  [15:0] result587;
wire  [15:0] result588;
wire  [15:0] result589;
wire  [15:0] result590;
wire  [15:0] result591;
wire  [15:0] result592;
wire  [15:0] result593;
wire  [15:0] result594;
wire  [15:0] result595;
wire  [15:0] result596;
wire  [15:0] result597;
wire  [15:0] result598;
wire  [15:0] result599;
wire  [15:0] result600;
wire  [15:0] result601;
wire  [15:0] result602;
wire  [15:0] result603;
wire  [15:0] result604;
wire  [15:0] result605;
wire  [15:0] result606;
wire  [15:0] result607;
wire  [15:0] result608;
wire  [15:0] result609;
wire  [15:0] result610;
wire  [15:0] result611;
wire  [15:0] result612;
wire  [15:0] result613;
wire  [15:0] result614;
wire  [15:0] result615;
wire  [15:0] result616;
wire  [15:0] result617;
wire  [15:0] result618;
wire  [15:0] result619;
wire  [15:0] result620;
wire  [15:0] result621;
wire  [15:0] result622;
wire  [15:0] result623;
wire  [15:0] result624;
wire  [15:0] result625;
wire  [15:0] result626;
wire  [15:0] result627;
wire  [15:0] result628;
wire  [15:0] result629;
wire  [15:0] result630;
wire  [15:0] result631;
wire  [15:0] result632;
wire  [15:0] result633;
wire  [15:0] result634;
wire  [15:0] result635;
wire  [15:0] result636;
wire  [15:0] result637;
wire  [15:0] result638;
wire  [15:0] result639;
wire  [15:0] result640;
wire  [15:0] result641;
wire  [15:0] result642;
wire  [15:0] result643;
wire  [15:0] result644;
wire  [15:0] result645;
wire  [15:0] result646;
wire  [15:0] result647;
wire  [15:0] result648;
wire  [15:0] result649;
wire  [15:0] result650;
wire  [15:0] result651;
wire  [15:0] result652;
wire  [15:0] result653;
wire  [15:0] result654;
wire  [15:0] result655;
wire  [15:0] result656;
wire  [15:0] result657;
wire  [15:0] result658;
wire  [15:0] result659;
wire  [15:0] result660;
wire  [15:0] result661;
wire  [15:0] result662;
wire  [15:0] result663;
wire  [15:0] result664;
wire  [15:0] result665;
wire  [15:0] result666;
wire  [15:0] result667;
wire  [15:0] result668;
wire  [15:0] result669;
wire  [15:0] result670;
wire  [15:0] result671;
wire  [15:0] result672;
wire  [15:0] result673;
wire  [15:0] result674;
wire  [15:0] result675;
wire  [15:0] result676;
wire  [15:0] result677;
wire  [15:0] result678;
wire  [15:0] result679;
wire  [15:0] result680;
wire  [15:0] result681;
wire  [15:0] result682;
wire  [15:0] result683;
wire  [15:0] result684;
wire  [15:0] result685;
wire  [15:0] result686;
wire  [15:0] result687;
wire  [15:0] result688;
wire  [15:0] result689;
wire  [15:0] result690;
wire  [15:0] result691;
wire  [15:0] result692;
wire  [15:0] result693;
wire  [15:0] result694;
wire  [15:0] result695;
wire  [15:0] result696;
wire  [15:0] result697;
wire  [15:0] result698;
wire  [15:0] result699;
wire  [15:0] result700;
wire  [15:0] result701;
wire  [15:0] result702;
wire  [15:0] result703;
wire  [15:0] result704;
wire  [15:0] result705;
wire  [15:0] result706;
wire  [15:0] result707;
wire  [15:0] result708;
wire  [15:0] result709;
wire  [15:0] result710;
wire  [15:0] result711;
wire  [15:0] result712;
wire  [15:0] result713;
wire  [15:0] result714;
wire  [15:0] result715;
wire  [15:0] result716;
wire  [15:0] result717;
wire  [15:0] result718;
wire  [15:0] result719;
wire  [15:0] result720;
wire  [15:0] result721;
wire  [15:0] result722;
wire  [15:0] result723;
wire  [15:0] result724;
wire  [15:0] result725;
wire  [15:0] result726;
wire  [15:0] result727;
wire  [15:0] result728;
wire  [15:0] result729;
wire  [15:0] result730;
wire  [15:0] result731;
wire  [15:0] result732;
wire  [15:0] result733;
wire  [15:0] result734;
wire  [15:0] result735;
wire  [15:0] result736;
wire  [15:0] result737;
wire  [15:0] result738;
wire  [15:0] result739;
wire  [15:0] result740;
wire  [15:0] result741;
wire  [15:0] result742;
wire  [15:0] result743;
wire  [15:0] result744;
wire  [15:0] result745;
wire  [15:0] result746;
wire  [15:0] result747;
wire  [15:0] result748;
wire  [15:0] result749;
wire  [15:0] result750;
wire  [15:0] result751;
wire  [15:0] result752;
wire  [15:0] result753;
wire  [15:0] result754;
wire  [15:0] result755;
wire  [15:0] result756;
wire  [15:0] result757;
wire  [15:0] result758;
wire  [15:0] result759;
wire  [15:0] result760;
wire  [15:0] result761;
wire  [15:0] result762;
wire  [15:0] result763;
wire  [15:0] result764;
wire  [15:0] result765;
wire  [15:0] result766;
wire  [15:0] result767;
wire  [15:0] result768;
wire  [15:0] result769;
wire  [15:0] result770;
wire  [15:0] result771;
wire  [15:0] result772;
wire  [15:0] result773;
wire  [15:0] result774;
wire  [15:0] result775;
wire  [15:0] result776;
wire  [15:0] result777;
wire  [15:0] result778;
wire  [15:0] result779;
wire  [15:0] result780;
wire  [15:0] result781;
wire  [15:0] result782;
wire  [15:0] result783;
wire  [15:0] result784;
wire  [15:0] result785;
wire  [15:0] result786;
wire  [15:0] result787;
wire  [15:0] result788;
wire  [15:0] result789;
wire  [15:0] result790;
wire  [15:0] result791;
wire  [15:0] result792;
wire  [15:0] result793;
wire  [15:0] result794;
wire  [15:0] result795;
wire  [15:0] result796;
wire  [15:0] result797;
wire  [15:0] result798;
wire  [15:0] result799;
wire  [15:0] result800;
wire  [15:0] result801;
wire  [15:0] result802;
wire  [15:0] result803;
wire  [15:0] result804;
wire  [15:0] result805;
wire  [15:0] result806;
wire  [15:0] result807;
wire  [15:0] result808;
wire  [15:0] result809;
wire  [15:0] result810;
wire  [15:0] result811;
wire  [15:0] result812;
wire  [15:0] result813;
wire  [15:0] result814;
wire  [15:0] result815;
wire  [15:0] result816;
wire  [15:0] result817;
wire  [15:0] result818;
wire  [15:0] result819;
wire  [15:0] result820;
wire  [15:0] result821;
wire  [15:0] result822;
wire  [15:0] result823;
wire  [15:0] result824;
wire  [15:0] result825;
wire  [15:0] result826;
wire  [15:0] result827;
wire  [15:0] result828;
wire  [15:0] result829;
wire  [15:0] result830;
wire  [15:0] result831;
wire  [15:0] result832;
wire  [15:0] result833;
wire  [15:0] result834;
wire  [15:0] result835;
wire  [15:0] result836;
wire  [15:0] result837;
wire  [15:0] result838;
wire  [15:0] result839;
wire  [15:0] result840;
wire  [15:0] result841;
wire  [15:0] result842;
wire  [15:0] result843;
wire  [15:0] result844;
wire  [15:0] result845;
wire  [15:0] result846;
wire  [15:0] result847;
wire  [15:0] result848;
wire  [15:0] result849;
wire  [15:0] result850;
wire  [15:0] result851;
wire  [15:0] result852;
wire  [15:0] result853;
wire  [15:0] result854;
wire  [15:0] result855;
wire  [15:0] result856;
wire  [15:0] result857;
wire  [15:0] result858;
wire  [15:0] result859;
wire  [15:0] result860;
wire  [15:0] result861;
wire  [15:0] result862;
wire  [15:0] result863;
wire  [15:0] result864;
wire  [15:0] result865;
wire  [15:0] result866;
wire  [15:0] result867;
wire  [15:0] result868;
wire  [15:0] result869;
wire  [15:0] result870;
wire  [15:0] result871;
wire  [15:0] result872;
wire  [15:0] result873;
wire  [15:0] result874;
wire  [15:0] result875;
wire  [15:0] result876;
wire  [15:0] result877;
wire  [15:0] result878;
wire  [15:0] result879;
wire  [15:0] result880;
wire  [15:0] result881;
wire  [15:0] result882;
wire  [15:0] result883;
wire  [15:0] result884;
wire  [15:0] result885;
wire  [15:0] result886;
wire  [15:0] result887;
wire  [15:0] result888;
wire  [15:0] result889;
wire  [15:0] result890;
wire  [15:0] result891;
wire  [15:0] result892;
wire  [15:0] result893;
wire  [15:0] result894;
wire  [15:0] result895;
wire  [15:0] result896;
wire  [15:0] result897;
wire  [15:0] result898;
wire  [15:0] result899;
wire  [15:0] result900;
wire  [15:0] result901;
wire  [15:0] result902;
wire  [15:0] result903;
wire  [15:0] result904;
wire  [15:0] result905;
wire  [15:0] result906;
wire  [15:0] result907;
wire  [15:0] result908;
wire  [15:0] result909;
wire  [15:0] result910;
wire  [15:0] result911;
wire  [15:0] result912;
wire  [15:0] result913;
wire  [15:0] result914;
wire  [15:0] result915;
wire  [15:0] result916;
wire  [15:0] result917;
wire  [15:0] result918;
wire  [15:0] result919;
wire  [15:0] result920;
wire  [15:0] result921;
wire  [15:0] result922;
wire  [15:0] result923;
wire  [15:0] result924;
wire  [15:0] result925;
wire  [15:0] result926;
wire  [15:0] result927;
wire  [15:0] result928;
wire  [15:0] result929;
wire  [15:0] result930;
wire  [15:0] result931;
wire  [15:0] result932;
wire  [15:0] result933;
wire  [15:0] result934;
wire  [15:0] result935;
wire  [15:0] result936;
wire  [15:0] result937;
wire  [15:0] result938;
wire  [15:0] result939;
wire  [15:0] result940;
wire  [15:0] result941;
wire  [15:0] result942;
wire  [15:0] result943;
wire  [15:0] result944;
wire  [15:0] result945;
wire  [15:0] result946;
wire  [15:0] result947;
wire  [15:0] result948;
wire  [15:0] result949;
wire  [15:0] result950;
wire  [15:0] result951;
wire  [15:0] result952;
wire  [15:0] result953;
wire  [15:0] result954;
wire  [15:0] result955;
wire  [15:0] result956;
wire  [15:0] result957;
wire  [15:0] result958;
wire  [15:0] result959;
wire  [15:0] result960;
wire  [15:0] result961;
wire  [15:0] result962;
wire  [15:0] result963;
wire  [15:0] result964;
wire  [15:0] result965;
wire  [15:0] result966;
wire  [15:0] result967;
wire  [15:0] result968;
wire  [15:0] result969;
wire  [15:0] result970;
wire  [15:0] result971;
wire  [15:0] result972;
wire  [15:0] result973;
wire  [15:0] result974;
wire  [15:0] result975;
wire  [15:0] result976;
wire  [15:0] result977;
wire  [15:0] result978;
wire  [15:0] result979;
wire  [15:0] result980;
wire  [15:0] result981;
wire  [15:0] result982;
wire  [15:0] result983;
wire  [15:0] result984;
wire  [15:0] result985;
wire  [15:0] result986;
wire  [15:0] result987;
wire  [15:0] result988;
wire  [15:0] result989;
wire  [15:0] result990;
wire  [15:0] result991;
wire  [15:0] result992;
wire  [15:0] result993;
wire  [15:0] result994;
wire  [15:0] result995;
wire  [15:0] result996;
wire  [15:0] result997;
wire  [15:0] result998;
wire  [15:0] result999;
wire  [15:0] result1000;
wire  [15:0] result1001;
wire  [15:0] result1002;
wire  [15:0] result1003;
wire  [15:0] result1004;
wire  [15:0] result1005;
wire  [15:0] result1006;
wire  [15:0] result1007;
wire  [15:0] result1008;
wire  [15:0] result1009;
wire  [15:0] result1010;
wire  [15:0] result1011;
wire  [15:0] result1012;
wire  [15:0] result1013;
wire  [15:0] result1014;
wire  [15:0] result1015;
wire  [15:0] result1016;
wire  [15:0] result1017;
wire  [15:0] result1018;
wire  [15:0] result1019;
wire  [15:0] result1020;
wire  [15:0] result1021;
wire  [15:0] result1022;
wire  [15:0] result1023;
wire  [15:0] result1024;
wire  [15:0] result1025;
wire  [15:0] result1026;
wire  [15:0] result1027;
wire  [15:0] result1028;
wire  [15:0] result1029;
wire  [15:0] result1030;
wire  [15:0] result1031;
wire  [15:0] result1032;
wire  [15:0] result1033;
wire  [15:0] result1034;
wire  [15:0] result1035;
wire  [15:0] result1036;
wire  [15:0] result1037;
wire  [15:0] result1038;
wire  [15:0] result1039;
wire  [15:0] result1040;
wire  [15:0] result1041;
wire  [15:0] result1042;
wire  [15:0] result1043;
wire  [15:0] result1044;
wire  [15:0] result1045;
wire  [15:0] result1046;
wire  [15:0] result1047;
wire  [15:0] result1048;
wire  [15:0] result1049;
wire  [15:0] result1050;
wire  [15:0] result1051;
wire  [15:0] result1052;
wire  [15:0] result1053;
wire  [15:0] result1054;
wire  [15:0] result1055;
wire  [15:0] result1056;
wire  [15:0] result1057;
wire  [15:0] result1058;
wire  [15:0] result1059;
wire  [15:0] result1060;
wire  [15:0] result1061;
wire  [15:0] result1062;
wire  [15:0] result1063;
wire  [15:0] result1064;
wire  [15:0] result1065;
wire  [15:0] result1066;
wire  [15:0] result1067;
wire  [15:0] result1068;
wire  [15:0] result1069;
wire  [15:0] result1070;
wire  [15:0] result1071;
wire  [15:0] result1072;
wire  [15:0] result1073;
wire  [15:0] result1074;
wire  [15:0] result1075;
wire  [15:0] result1076;
wire  [15:0] result1077;
wire  [15:0] result1078;
wire  [15:0] result1079;
wire  [15:0] result1080;
wire  [15:0] result1081;
wire  [15:0] result1082;
wire  [15:0] result1083;
wire  [15:0] result1084;
wire  [15:0] result1085;
wire  [15:0] result1086;
wire  [15:0] result1087;
wire  [15:0] result1088;
wire  [15:0] result1089;
wire  [15:0] result1090;
wire  [15:0] result1091;
wire  [15:0] result1092;
wire  [15:0] result1093;
wire  [15:0] result1094;
wire  [15:0] result1095;
wire  [15:0] result1096;
wire  [15:0] result1097;
wire  [15:0] result1098;
wire  [15:0] result1099;
wire  [15:0] result1100;
wire  [15:0] result1101;
wire  [15:0] result1102;
wire  [15:0] result1103;
wire  [15:0] result1104;
wire  [15:0] result1105;
wire  [15:0] result1106;
wire  [15:0] result1107;
wire  [15:0] result1108;
wire  [15:0] result1109;
wire  [15:0] result1110;
wire  [15:0] result1111;
wire  [15:0] result1112;
wire  [15:0] result1113;
wire  [15:0] result1114;
wire  [15:0] result1115;
wire  [15:0] result1116;
wire  [15:0] result1117;
wire  [15:0] result1118;
wire  [15:0] result1119;
wire  [15:0] result1120;
wire  [15:0] result1121;
wire  [15:0] result1122;
wire  [15:0] result1123;
wire  [15:0] result1124;
wire  [15:0] result1125;
wire  [15:0] result1126;
wire  [15:0] result1127;
wire  [15:0] result1128;
wire  [15:0] result1129;
wire  [15:0] result1130;
wire  [15:0] result1131;
wire  [15:0] result1132;
wire  [15:0] result1133;
wire  [15:0] result1134;
wire  [15:0] result1135;
wire  [15:0] result1136;
wire  [15:0] result1137;
wire  [15:0] result1138;
wire  [15:0] result1139;
wire  [15:0] result1140;
wire  [15:0] result1141;
wire  [15:0] result1142;
wire  [15:0] result1143;
wire  [15:0] result1144;
wire  [15:0] result1145;
wire  [15:0] result1146;
wire  [15:0] result1147;
wire  [15:0] result1148;
wire  [15:0] result1149;
wire  [15:0] result1150;
wire  [15:0] result1151;
wire  [15:0] result1152;
wire  [15:0] result1153;
wire  [15:0] result1154;
wire  [15:0] result1155;
wire  [15:0] result1156;
wire  [15:0] result1157;
wire  [15:0] result1158;
wire  [15:0] result1159;
wire  [15:0] result1160;
wire  [15:0] result1161;
wire  [15:0] result1162;
wire  [15:0] result1163;
wire  [15:0] result1164;
wire  [15:0] result1165;
wire  [15:0] result1166;
wire  [15:0] result1167;
wire  [15:0] result1168;
wire  [15:0] result1169;
wire  [15:0] result1170;
wire  [15:0] result1171;
wire  [15:0] result1172;
wire  [15:0] result1173;
wire  [15:0] result1174;
wire  [15:0] result1175;
wire  [15:0] result1176;
wire  [15:0] result1177;
wire  [15:0] result1178;
wire  [15:0] result1179;
wire  [15:0] result1180;
wire  [15:0] result1181;
wire  [15:0] result1182;
wire  [15:0] result1183;
wire  [15:0] result1184;
wire  [15:0] result1185;
wire  [15:0] result1186;
wire  [15:0] result1187;
wire  [15:0] result1188;
wire  [15:0] result1189;
wire  [15:0] result1190;
wire  [15:0] result1191;
wire  [15:0] result1192;
wire  [15:0] result1193;
wire  [15:0] result1194;
wire  [15:0] result1195;
wire  [15:0] result1196;
wire  [15:0] result1197;
wire  [15:0] result1198;
wire  [15:0] result1199;
wire  [15:0] result1200;
wire  [15:0] result1201;
wire  [15:0] result1202;
wire  [15:0] result1203;
wire  [15:0] result1204;
wire  [15:0] result1205;
wire  [15:0] result1206;
wire  [15:0] result1207;
wire  [15:0] result1208;
wire  [15:0] result1209;
wire  [15:0] result1210;
wire  [15:0] result1211;
wire  [15:0] result1212;
wire  [15:0] result1213;
wire  [15:0] result1214;
wire  [15:0] result1215;
wire  [15:0] result1216;
wire  [15:0] result1217;
wire  [15:0] result1218;
wire  [15:0] result1219;
wire  [15:0] result1220;
wire  [15:0] result1221;
wire  [15:0] result1222;
wire  [15:0] result1223;
wire  [15:0] result1224;
wire  [15:0] result1225;
wire  [15:0] result1226;
wire  [15:0] result1227;
wire  [15:0] result1228;
wire  [15:0] result1229;
wire  [15:0] result1230;
wire  [15:0] result1231;
wire  [15:0] result1232;
wire  [15:0] result1233;
wire  [15:0] result1234;
wire  [15:0] result1235;
wire  [15:0] result1236;
wire  [15:0] result1237;
wire  [15:0] result1238;
wire  [15:0] result1239;
wire  [15:0] result1240;
wire  [15:0] result1241;
wire  [15:0] result1242;
wire  [15:0] result1243;
wire  [15:0] result1244;
wire  [15:0] result1245;
wire  [15:0] result1246;
wire  [15:0] result1247;
wire  [15:0] result1248;
wire  [15:0] result1249;
wire  [15:0] result1250;
wire  [15:0] result1251;
wire  [15:0] result1252;
wire  [15:0] result1253;
wire  [15:0] result1254;
wire  [15:0] result1255;
wire  [15:0] result1256;
wire  [15:0] result1257;
wire  [15:0] result1258;
wire  [15:0] result1259;
wire  [15:0] result1260;
wire  [15:0] result1261;
wire  [15:0] result1262;
wire  [15:0] result1263;
wire  [15:0] result1264;
wire  [15:0] result1265;
wire  [15:0] result1266;
wire  [15:0] result1267;
wire  [15:0] result1268;
wire  [15:0] result1269;
wire  [15:0] result1270;
wire  [15:0] result1271;
wire  [15:0] result1272;
wire  [15:0] result1273;
wire  [15:0] result1274;
wire  [15:0] result1275;
wire  [15:0] result1276;
wire  [15:0] result1277;
wire  [15:0] result1278;
wire  [15:0] result1279;
wire  [15:0] result1280;
wire  [15:0] result1281;
wire  [15:0] result1282;
wire  [15:0] result1283;
wire  [15:0] result1284;
wire  [15:0] result1285;
wire  [15:0] result1286;
wire  [15:0] result1287;
wire  [15:0] result1288;
wire  [15:0] result1289;
wire  [15:0] result1290;
wire  [15:0] result1291;
wire  [15:0] result1292;
wire  [15:0] result1293;
wire  [15:0] result1294;
wire  [15:0] result1295;
wire  [15:0] result1296;
wire  [15:0] result1297;
wire  [15:0] result1298;
wire  [15:0] result1299;
wire  [15:0] result1300;
wire  [15:0] result1301;
wire  [15:0] result1302;
wire  [15:0] result1303;
wire  [15:0] result1304;
wire  [15:0] result1305;
wire  [15:0] result1306;
wire  [15:0] result1307;
wire  [15:0] result1308;
wire  [15:0] result1309;
wire  [15:0] result1310;
wire  [15:0] result1311;
wire  [15:0] result1312;
wire  [15:0] result1313;
wire  [15:0] result1314;
wire  [15:0] result1315;
wire  [15:0] result1316;
wire  [15:0] result1317;
wire  [15:0] result1318;
wire  [15:0] result1319;
wire  [15:0] result1320;
wire  [15:0] result1321;
wire  [15:0] result1322;
wire  [15:0] result1323;
wire  [15:0] result1324;
wire  [15:0] result1325;
wire  [15:0] result1326;
wire  [15:0] result1327;
wire  [15:0] result1328;
wire  [15:0] result1329;
wire  [15:0] result1330;
wire  [15:0] result1331;
wire  [15:0] result1332;
wire  [15:0] result1333;
wire  [15:0] result1334;
wire  [15:0] result1335;
wire  [15:0] result1336;
wire  [15:0] result1337;
wire  [15:0] result1338;
wire  [15:0] result1339;
wire  [15:0] result1340;
wire  [15:0] result1341;
wire  [15:0] result1342;
wire  [15:0] result1343;
wire  [15:0] result1344;
wire  [15:0] result1345;
wire  [15:0] result1346;
wire  [15:0] result1347;
wire  [15:0] result1348;
wire  [15:0] result1349;
wire  [15:0] result1350;
wire  [15:0] result1351;
wire  [15:0] result1352;
wire  [15:0] result1353;
wire  [15:0] result1354;
wire  [15:0] result1355;
wire  [15:0] result1356;
wire  [15:0] result1357;
wire  [15:0] result1358;
wire  [15:0] result1359;
wire  [15:0] result1360;
wire  [15:0] result1361;
wire  [15:0] result1362;
wire  [15:0] result1363;
wire  [15:0] result1364;
wire  [15:0] result1365;
wire  [15:0] result1366;
wire  [15:0] result1367;
wire  [15:0] result1368;
wire  [15:0] result1369;
wire  [15:0] result1370;
wire  [15:0] result1371;
wire  [15:0] result1372;
wire  [15:0] result1373;
wire  [15:0] result1374;
wire  [15:0] result1375;
wire  [15:0] result1376;
wire  [15:0] result1377;
wire  [15:0] result1378;
wire  [15:0] result1379;
wire  [15:0] result1380;
wire  [15:0] result1381;
wire  [15:0] result1382;
wire  [15:0] result1383;
wire  [15:0] result1384;
wire  [15:0] result1385;
wire  [15:0] result1386;
wire  [15:0] result1387;
wire  [15:0] result1388;
wire  [15:0] result1389;
wire  [15:0] result1390;
wire  [15:0] result1391;
wire  [15:0] result1392;
wire  [15:0] result1393;
wire  [15:0] result1394;
wire  [15:0] result1395;
wire  [15:0] result1396;
wire  [15:0] result1397;
wire  [15:0] result1398;
wire  [15:0] result1399;
wire  [15:0] result1400;
wire  [15:0] result1401;
wire  [15:0] result1402;
wire  [15:0] result1403;
wire  [15:0] result1404;
wire  [15:0] result1405;
wire  [15:0] result1406;
wire  [15:0] result1407;
wire  [15:0] result1408;
wire  [15:0] result1409;
wire  [15:0] result1410;
wire  [15:0] result1411;
wire  [15:0] result1412;
wire  [15:0] result1413;
wire  [15:0] result1414;
wire  [15:0] result1415;
wire  [15:0] result1416;
wire  [15:0] result1417;
wire  [15:0] result1418;
wire  [15:0] result1419;
wire  [15:0] result1420;
wire  [15:0] result1421;
wire  [15:0] result1422;
wire  [15:0] result1423;
wire  [15:0] result1424;
wire  [15:0] result1425;
wire  [15:0] result1426;
wire  [15:0] result1427;
wire  [15:0] result1428;
wire  [15:0] result1429;
wire  [15:0] result1430;
wire  [15:0] result1431;
wire  [15:0] result1432;
wire  [15:0] result1433;
wire  [15:0] result1434;
wire  [15:0] result1435;
wire  [15:0] result1436;
wire  [15:0] result1437;
wire  [15:0] result1438;
wire  [15:0] result1439;
wire  [15:0] result1440;
wire  [15:0] result1441;
wire  [15:0] result1442;
wire  [15:0] result1443;
wire  [15:0] result1444;
wire  [15:0] result1445;
wire  [15:0] result1446;
wire  [15:0] result1447;
wire  [15:0] result1448;
wire  [15:0] result1449;
wire  [15:0] result1450;
wire  [15:0] result1451;
wire  [15:0] result1452;
wire  [15:0] result1453;
wire  [15:0] result1454;
wire  [15:0] result1455;
wire  [15:0] result1456;
wire  [15:0] result1457;
wire  [15:0] result1458;
wire  [15:0] result1459;
wire  [15:0] result1460;
wire  [15:0] result1461;
wire  [15:0] result1462;
wire  [15:0] result1463;
wire  [15:0] result1464;
wire  [15:0] result1465;
wire  [15:0] result1466;
wire  [15:0] result1467;
wire  [15:0] result1468;
wire  [15:0] result1469;
wire  [15:0] result1470;
wire  [15:0] result1471;
wire  [15:0] result1472;
wire  [15:0] result1473;
wire  [15:0] result1474;
wire  [15:0] result1475;
wire  [15:0] result1476;
wire  [15:0] result1477;
wire  [15:0] result1478;
wire  [15:0] result1479;
wire  [15:0] result1480;
wire  [15:0] result1481;
wire  [15:0] result1482;
wire  [15:0] result1483;
wire  [15:0] result1484;
wire  [15:0] result1485;
wire  [15:0] result1486;
wire  [15:0] result1487;
wire  [15:0] result1488;
wire  [15:0] result1489;
wire  [15:0] result1490;
wire  [15:0] result1491;
wire  [15:0] result1492;
wire  [15:0] result1493;
wire  [15:0] result1494;
wire  [15:0] result1495;
wire  [15:0] result1496;
wire  [15:0] result1497;
wire  [15:0] result1498;
wire  [15:0] result1499;
wire  [15:0] result1500;
wire  [15:0] result1501;
wire  [15:0] result1502;
wire  [15:0] result1503;
wire  [15:0] result1504;
wire  [15:0] result1505;
wire  [15:0] result1506;
wire  [15:0] result1507;
wire  [15:0] result1508;
wire  [15:0] result1509;
wire  [15:0] result1510;
wire  [15:0] result1511;
wire  [15:0] result1512;
wire  [15:0] result1513;
wire  [15:0] result1514;
wire  [15:0] result1515;
wire  [15:0] result1516;
wire  [15:0] result1517;
wire  [15:0] result1518;
wire  [15:0] result1519;
wire  [15:0] result1520;
wire  [15:0] result1521;
wire  [15:0] result1522;
wire  [15:0] result1523;
wire  [15:0] result1524;
wire  [15:0] result1525;
wire  [15:0] result1526;
wire  [15:0] result1527;
wire  [15:0] result1528;
wire  [15:0] result1529;
wire  [15:0] result1530;
wire  [15:0] result1531;
wire  [15:0] result1532;
wire  [15:0] result1533;
wire  [15:0] result1534;
wire  [15:0] result1535;
wire  [15:0] result1536;
wire  [15:0] result1537;
wire  [15:0] result1538;
wire  [15:0] result1539;
wire  [15:0] result1540;
wire  [15:0] result1541;
wire  [15:0] result1542;
wire  [15:0] result1543;
wire  [15:0] result1544;
wire  [15:0] result1545;
wire  [15:0] result1546;
wire  [15:0] result1547;
wire  [15:0] result1548;
wire  [15:0] result1549;
wire  [15:0] result1550;
wire  [15:0] result1551;
wire  [15:0] result1552;
wire  [15:0] result1553;
wire  [15:0] result1554;
wire  [15:0] result1555;
wire  [15:0] result1556;
wire  [15:0] result1557;
wire  [15:0] result1558;
wire  [15:0] result1559;
wire  [15:0] result1560;
wire  [15:0] result1561;
wire  [15:0] result1562;
wire  [15:0] result1563;
wire  [15:0] result1564;
wire  [15:0] result1565;
wire  [15:0] result1566;
wire  [15:0] result1567;
wire  [15:0] result1568;
wire  [15:0] result1569;
wire  [15:0] result1570;
wire  [15:0] result1571;
wire  [15:0] result1572;
wire  [15:0] result1573;
wire  [15:0] result1574;
wire  [15:0] result1575;
wire  [15:0] result1576;
wire  [15:0] result1577;
wire  [15:0] result1578;
wire  [15:0] result1579;
wire  [15:0] result1580;
wire  [15:0] result1581;
wire  [15:0] result1582;
wire  [15:0] result1583;
wire  [15:0] result1584;
wire  [15:0] result1585;
wire  [15:0] result1586;
wire  [15:0] result1587;
wire  [15:0] result1588;
wire  [15:0] result1589;
wire  [15:0] result1590;
wire  [15:0] result1591;
wire  [15:0] result1592;
wire  [15:0] result1593;
wire  [15:0] result1594;
wire  [15:0] result1595;
wire  [15:0] result1596;
wire  [15:0] result1597;
wire  [15:0] result1598;
wire  [15:0] result1599;
wire  [15:0] result1600;
wire  [15:0] result1601;
wire  [15:0] result1602;
wire  [15:0] result1603;
wire  [15:0] result1604;
wire  [15:0] result1605;
wire  [15:0] result1606;
wire  [15:0] result1607;
wire  [15:0] result1608;
wire  [15:0] result1609;
wire  [15:0] result1610;
wire  [15:0] result1611;
wire  [15:0] result1612;
wire  [15:0] result1613;
wire  [15:0] result1614;
wire  [15:0] result1615;
wire  [15:0] result1616;
wire  [15:0] result1617;
wire  [15:0] result1618;
wire  [15:0] result1619;
wire  [15:0] result1620;
wire  [15:0] result1621;
wire  [15:0] result1622;
wire  [15:0] result1623;
wire  [15:0] result1624;
wire  [15:0] result1625;
wire  [15:0] result1626;
wire  [15:0] result1627;
wire  [15:0] result1628;
wire  [15:0] result1629;
wire  [15:0] result1630;
wire  [15:0] result1631;
wire  [15:0] result1632;
wire  [15:0] result1633;
wire  [15:0] result1634;
wire  [15:0] result1635;
wire  [15:0] result1636;
wire  [15:0] result1637;
wire  [15:0] result1638;
wire  [15:0] result1639;
wire  [15:0] result1640;
wire  [15:0] result1641;
wire  [15:0] result1642;
wire  [15:0] result1643;
wire  [15:0] result1644;
wire  [15:0] result1645;
wire  [15:0] result1646;
wire  [15:0] result1647;
wire  [15:0] result1648;
wire  [15:0] result1649;
wire  [15:0] result1650;
wire  [15:0] result1651;
wire  [15:0] result1652;
wire  [15:0] result1653;
wire  [15:0] result1654;
wire  [15:0] result1655;
wire  [15:0] result1656;
wire  [15:0] result1657;
wire  [15:0] result1658;
wire  [15:0] result1659;
wire  [15:0] result1660;
wire  [15:0] result1661;
wire  [15:0] result1662;
wire  [15:0] result1663;
wire  [15:0] result1664;
wire  [15:0] result1665;
wire  [15:0] result1666;
wire  [15:0] result1667;
wire  [15:0] result1668;
wire  [15:0] result1669;
wire  [15:0] result1670;
wire  [15:0] result1671;
wire  [15:0] result1672;
wire  [15:0] result1673;
wire  [15:0] result1674;
wire  [15:0] result1675;
wire  [15:0] result1676;
wire  [15:0] result1677;
wire  [15:0] result1678;
wire  [15:0] result1679;
wire  [15:0] result1680;
wire  [15:0] result1681;
wire  [15:0] result1682;
wire  [15:0] result1683;
wire  [15:0] result1684;
wire  [15:0] result1685;
wire  [15:0] result1686;
wire  [15:0] result1687;
wire  [15:0] result1688;
wire  [15:0] result1689;
wire  [15:0] result1690;
wire  [15:0] result1691;
wire  [15:0] result1692;
wire  [15:0] result1693;
wire  [15:0] result1694;
wire  [15:0] result1695;
wire  [15:0] result1696;
wire  [15:0] result1697;
wire  [15:0] result1698;
wire  [15:0] result1699;
wire  [15:0] result1700;
wire  [15:0] result1701;
wire  [15:0] result1702;
wire  [15:0] result1703;
wire  [15:0] result1704;
wire  [15:0] result1705;
wire  [15:0] result1706;
wire  [15:0] result1707;
wire  [15:0] result1708;
wire  [15:0] result1709;
wire  [15:0] result1710;
wire  [15:0] result1711;
wire  [15:0] result1712;
wire  [15:0] result1713;
wire  [15:0] result1714;
wire  [15:0] result1715;
wire  [15:0] result1716;
wire  [15:0] result1717;
wire  [15:0] result1718;
wire  [15:0] result1719;
wire  [15:0] result1720;
wire  [15:0] result1721;
wire  [15:0] result1722;
wire  [15:0] result1723;
wire  [15:0] result1724;
wire  [15:0] result1725;
wire  [15:0] result1726;
wire  [15:0] result1727;
wire  [15:0] result1728;
wire  [15:0] result1729;
wire  [15:0] result1730;
wire  [15:0] result1731;
wire  [15:0] result1732;
wire  [15:0] result1733;
wire  [15:0] result1734;
wire  [15:0] result1735;
wire  [15:0] result1736;
wire  [15:0] result1737;
wire  [15:0] result1738;
wire  [15:0] result1739;
wire  [15:0] result1740;
wire  [15:0] result1741;
wire  [15:0] result1742;
wire  [15:0] result1743;
wire  [15:0] result1744;
wire  [15:0] result1745;
wire  [15:0] result1746;
wire  [15:0] result1747;
wire  [15:0] result1748;
wire  [15:0] result1749;
wire  [15:0] result1750;
wire  [15:0] result1751;
wire  [15:0] result1752;
wire  [15:0] result1753;
wire  [15:0] result1754;
wire  [15:0] result1755;
wire  [15:0] result1756;
wire  [15:0] result1757;
wire  [15:0] result1758;
wire  [15:0] result1759;
wire  [15:0] result1760;
wire  [15:0] result1761;
wire  [15:0] result1762;
wire  [15:0] result1763;
wire  [15:0] result1764;
wire  [15:0] result1765;
wire  [15:0] result1766;
wire  [15:0] result1767;
wire  [15:0] result1768;
wire  [15:0] result1769;
wire  [15:0] result1770;
wire  [15:0] result1771;
wire  [15:0] result1772;
wire  [15:0] result1773;
wire  [15:0] result1774;
wire  [15:0] result1775;
wire  [15:0] result1776;
wire  [15:0] result1777;
wire  [15:0] result1778;
wire  [15:0] result1779;
wire  [15:0] result1780;
wire  [15:0] result1781;
wire  [15:0] result1782;
wire  [15:0] result1783;
wire  [15:0] result1784;
wire  [15:0] result1785;
wire  [15:0] result1786;
wire  [15:0] result1787;
wire  [15:0] result1788;
wire  [15:0] result1789;
wire  [15:0] result1790;
wire  [15:0] result1791;
wire  [15:0] result1792;
wire  [15:0] result1793;
wire  [15:0] result1794;
wire  [15:0] result1795;
wire  [15:0] result1796;
wire  [15:0] result1797;
wire  [15:0] result1798;
wire  [15:0] result1799;
wire  [15:0] result1800;
wire  [15:0] result1801;
wire  [15:0] result1802;
wire  [15:0] result1803;
wire  [15:0] result1804;
wire  [15:0] result1805;
wire  [15:0] result1806;
wire  [15:0] result1807;
wire  [15:0] result1808;
wire  [15:0] result1809;
wire  [15:0] result1810;
wire  [15:0] result1811;
wire  [15:0] result1812;
wire  [15:0] result1813;
wire  [15:0] result1814;
wire  [15:0] result1815;
wire  [15:0] result1816;
wire  [15:0] result1817;
wire  [15:0] result1818;
wire  [15:0] result1819;
wire  [15:0] result1820;
wire  [15:0] result1821;
wire  [15:0] result1822;
wire  [15:0] result1823;
wire  [15:0] result1824;
wire  [15:0] result1825;
wire  [15:0] result1826;
wire  [15:0] result1827;
wire  [15:0] result1828;
wire  [15:0] result1829;
wire  [15:0] result1830;
wire  [15:0] result1831;
wire  [15:0] result1832;
wire  [15:0] result1833;
wire  [15:0] result1834;
wire  [15:0] result1835;
wire  [15:0] result1836;
wire  [15:0] result1837;
wire  [15:0] result1838;
wire  [15:0] result1839;
wire  [15:0] result1840;
wire  [15:0] result1841;
wire  [15:0] result1842;
wire  [15:0] result1843;
wire  [15:0] result1844;
wire  [15:0] result1845;
wire  [15:0] result1846;
wire  [15:0] result1847;
wire  [15:0] result1848;
wire  [15:0] result1849;
wire  [15:0] result1850;
wire  [15:0] result1851;
wire  [15:0] result1852;
wire  [15:0] result1853;
wire  [15:0] result1854;
wire  [15:0] result1855;
wire  [15:0] result1856;
wire  [15:0] result1857;
wire  [15:0] result1858;
wire  [15:0] result1859;
wire  [15:0] result1860;
wire  [15:0] result1861;
wire  [15:0] result1862;
wire  [15:0] result1863;
wire  [15:0] result1864;
wire  [15:0] result1865;
wire  [15:0] result1866;
wire  [15:0] result1867;
wire  [15:0] result1868;
wire  [15:0] result1869;
wire  [15:0] result1870;
wire  [15:0] result1871;
wire  [15:0] result1872;
wire  [15:0] result1873;
wire  [15:0] result1874;
wire  [15:0] result1875;
wire  [15:0] result1876;
wire  [15:0] result1877;
wire  [15:0] result1878;
wire  [15:0] result1879;
wire  [15:0] result1880;
wire  [15:0] result1881;
wire  [15:0] result1882;
wire  [15:0] result1883;
wire  [15:0] result1884;
wire  [15:0] result1885;
wire  [15:0] result1886;
wire  [15:0] result1887;
wire  [15:0] result1888;
wire  [15:0] result1889;
wire  [15:0] result1890;
wire  [15:0] result1891;
wire  [15:0] result1892;
wire  [15:0] result1893;
wire  [15:0] result1894;
wire  [15:0] result1895;
wire  [15:0] result1896;
wire  [15:0] result1897;
wire  [15:0] result1898;
wire  [15:0] result1899;
wire  [15:0] result1900;
wire  [15:0] result1901;
wire  [15:0] result1902;
wire  [15:0] result1903;
wire  [15:0] result1904;
wire  [15:0] result1905;
wire  [15:0] result1906;
wire  [15:0] result1907;
wire  [15:0] result1908;
wire  [15:0] result1909;
wire  [15:0] result1910;
wire  [15:0] result1911;
wire  [15:0] result1912;
wire  [15:0] result1913;
wire  [15:0] result1914;
wire  [15:0] result1915;
wire  [15:0] result1916;
wire  [15:0] result1917;
wire  [15:0] result1918;
wire  [15:0] result1919;
wire  [15:0] result1920;
wire  [15:0] result1921;
wire  [15:0] result1922;
wire  [15:0] result1923;
wire  [15:0] result1924;
wire  [15:0] result1925;
wire  [15:0] result1926;
wire  [15:0] result1927;
wire  [15:0] result1928;
wire  [15:0] result1929;
wire  [15:0] result1930;
wire  [15:0] result1931;
wire  [15:0] result1932;
wire  [15:0] result1933;
wire  [15:0] result1934;
wire  [15:0] result1935;
wire  [15:0] result1936;
wire  [15:0] result1937;
wire  [15:0] result1938;
wire  [15:0] result1939;
wire  [15:0] result1940;
wire  [15:0] result1941;
wire  [15:0] result1942;
wire  [15:0] result1943;
wire  [15:0] result1944;
wire  [15:0] result1945;
wire  [15:0] result1946;
wire  [15:0] result1947;
wire  [15:0] result1948;
wire  [15:0] result1949;
wire  [15:0] result1950;
wire  [15:0] result1951;
wire  [15:0] result1952;
wire  [15:0] result1953;
wire  [15:0] result1954;
wire  [15:0] result1955;
wire  [15:0] result1956;
wire  [15:0] result1957;
wire  [15:0] result1958;
wire  [15:0] result1959;
wire  [15:0] result1960;
wire  [15:0] result1961;
wire  [15:0] result1962;
wire  [15:0] result1963;
wire  [15:0] result1964;
wire  [15:0] result1965;
wire  [15:0] result1966;
wire  [15:0] result1967;
wire  [15:0] result1968;
wire  [15:0] result1969;
wire  [15:0] result1970;
wire  [15:0] result1971;
wire  [15:0] result1972;
wire  [15:0] result1973;
wire  [15:0] result1974;
wire  [15:0] result1975;
wire  [15:0] result1976;
wire  [15:0] result1977;
wire  [15:0] result1978;
wire  [15:0] result1979;
wire  [15:0] result1980;
wire  [15:0] result1981;
wire  [15:0] result1982;
wire  [15:0] result1983;
wire  [15:0] result1984;
wire  [15:0] result1985;
wire  [15:0] result1986;
wire  [15:0] result1987;
wire  [15:0] result1988;
wire  [15:0] result1989;
wire  [15:0] result1990;
wire  [15:0] result1991;
wire  [15:0] result1992;
wire  [15:0] result1993;
wire  [15:0] result1994;
wire  [15:0] result1995;
wire  [15:0] result1996;
wire  [15:0] result1997;
wire  [15:0] result1998;
wire  [15:0] result1999;
wire  [15:0] result2000;
wire  [15:0] result2001;
wire  [15:0] result2002;
wire  [15:0] result2003;
wire  [15:0] result2004;
wire  [15:0] result2005;
wire  [15:0] result2006;
wire  [15:0] result2007;
wire  [15:0] result2008;
wire  [15:0] result2009;
wire  [15:0] result2010;
wire  [15:0] result2011;
wire  [15:0] result2012;
wire  [15:0] result2013;
wire  [15:0] result2014;
wire  [15:0] result2015;
wire  [15:0] result2016;
wire  [15:0] result2017;
wire  [15:0] result2018;
wire  [15:0] result2019;
wire  [15:0] result2020;
wire  [15:0] result2021;
wire  [15:0] result2022;
wire  [15:0] result2023;
wire  [15:0] result2024;
wire  [15:0] result2025;
wire  [15:0] result2026;
wire  [15:0] result2027;
wire  [15:0] result2028;
wire  [15:0] result2029;
wire  [15:0] result2030;
wire  [15:0] result2031;
wire  [15:0] result2032;
wire  [15:0] result2033;
wire  [15:0] result2034;
wire  [15:0] result2035;
wire  [15:0] result2036;
wire  [15:0] result2037;
wire  [15:0] result2038;
wire  [15:0] result2039;
wire  [15:0] result2040;
wire  [15:0] result2041;
wire  [15:0] result2042;
wire  [15:0] result2043;
wire  [15:0] result2044;
wire  [15:0] result2045;
wire  [15:0] result2046;
wire  [15:0] result2047;
wire  [15:0] result2048;
wire  [15:0] result2049;
wire  [15:0] result2050;
wire  [15:0] result2051;
wire  [15:0] result2052;
wire  [15:0] result2053;
wire  [15:0] result2054;
wire  [15:0] result2055;
wire  [15:0] result2056;
wire  [15:0] result2057;
wire  [15:0] result2058;
wire  [15:0] result2059;
wire  [15:0] result2060;
wire  [15:0] result2061;
wire  [15:0] result2062;
wire  [15:0] result2063;
wire  [15:0] result2064;
wire  [15:0] result2065;
wire  [15:0] result2066;
wire  [15:0] result2067;
wire  [15:0] result2068;
wire  [15:0] result2069;
wire  [15:0] result2070;
wire  [15:0] result2071;
wire  [15:0] result2072;
wire  [15:0] result2073;
wire  [15:0] result2074;
wire  [15:0] result2075;
wire  [15:0] result2076;
wire  [15:0] result2077;
wire  [15:0] result2078;
wire  [15:0] result2079;
wire  [15:0] result2080;
wire  [15:0] result2081;
wire  [15:0] result2082;
wire  [15:0] result2083;
wire  [15:0] result2084;
wire  [15:0] result2085;
wire  [15:0] result2086;
wire  [15:0] result2087;
wire  [15:0] result2088;
wire  [15:0] result2089;
wire  [15:0] result2090;
wire  [15:0] result2091;
wire  [15:0] result2092;
wire  [15:0] result2093;
wire  [15:0] result2094;
wire  [15:0] result2095;
wire  [15:0] result2096;
wire  [15:0] result2097;
wire  [15:0] result2098;
wire  [15:0] result2099;
wire  [15:0] result2100;
wire  [15:0] result2101;
wire  [15:0] result2102;
wire  [15:0] result2103;
wire  [15:0] result2104;
wire  [15:0] result2105;
wire  [15:0] result2106;
wire  [15:0] result2107;
wire  [15:0] result2108;
wire  [15:0] result2109;
wire  [15:0] result2110;
wire  [15:0] result2111;
wire  [15:0] result2112;
wire  [15:0] result2113;
wire  [15:0] result2114;
wire  [15:0] result2115;
wire  [15:0] result2116;
wire  [15:0] result2117;
wire  [15:0] result2118;
wire  [15:0] result2119;
wire  [15:0] result2120;
wire  [15:0] result2121;
wire  [15:0] result2122;
wire  [15:0] result2123;
wire  [15:0] result2124;
wire  [15:0] result2125;
wire  [15:0] result2126;
wire  [15:0] result2127;
wire  [15:0] result2128;
wire  [15:0] result2129;
wire  [15:0] result2130;
wire  [15:0] result2131;
wire  [15:0] result2132;
wire  [15:0] result2133;
wire  [15:0] result2134;
wire  [15:0] result2135;
wire  [15:0] result2136;
wire  [15:0] result2137;
wire  [15:0] result2138;
wire  [15:0] result2139;
wire  [15:0] result2140;
wire  [15:0] result2141;
wire  [15:0] result2142;
wire  [15:0] result2143;
wire  [15:0] result2144;
wire  [15:0] result2145;
wire  [15:0] result2146;
wire  [15:0] result2147;
wire  [15:0] result2148;
wire  [15:0] result2149;
wire  [15:0] result2150;
wire  [15:0] result2151;
wire  [15:0] result2152;
wire  [15:0] result2153;
wire  [15:0] result2154;
wire  [15:0] result2155;
wire  [15:0] result2156;
wire  [15:0] result2157;
wire  [15:0] result2158;
wire  [15:0] result2159;
wire  [15:0] result2160;
wire  [15:0] result2161;
wire  [15:0] result2162;
wire  [15:0] result2163;
wire  [15:0] result2164;
wire  [15:0] result2165;
wire  [15:0] result2166;
wire  [15:0] result2167;
wire  [15:0] result2168;
wire  [15:0] result2169;
wire  [15:0] result2170;
wire  [15:0] result2171;
wire  [15:0] result2172;
wire  [15:0] result2173;
wire  [15:0] result2174;
wire  [15:0] result2175;
wire  [15:0] result2176;
wire  [15:0] result2177;
wire  [15:0] result2178;
wire  [15:0] result2179;
wire  [15:0] result2180;
wire  [15:0] result2181;
wire  [15:0] result2182;
wire  [15:0] result2183;
wire  [15:0] result2184;
wire  [15:0] result2185;
wire  [15:0] result2186;
wire  [15:0] result2187;
wire  [15:0] result2188;
wire  [15:0] result2189;
wire  [15:0] result2190;
wire  [15:0] result2191;
wire  [15:0] result2192;
wire  [15:0] result2193;
wire  [15:0] result2194;
wire  [15:0] result2195;
wire  [15:0] result2196;
wire  [15:0] result2197;
wire  [15:0] result2198;
wire  [15:0] result2199;
wire  [15:0] result2200;
wire  [15:0] result2201;
wire  [15:0] result2202;
wire  [15:0] result2203;
wire  [15:0] result2204;
wire  [15:0] result2205;
wire  [15:0] result2206;
wire  [15:0] result2207;
wire  [15:0] result2208;
wire  [15:0] result2209;
wire  [15:0] result2210;
wire  [15:0] result2211;
wire  [15:0] result2212;
wire  [15:0] result2213;
wire  [15:0] result2214;
wire  [15:0] result2215;
wire  [15:0] result2216;
wire  [15:0] result2217;
wire  [15:0] result2218;
wire  [15:0] result2219;
wire  [15:0] result2220;
wire  [15:0] result2221;
wire  [15:0] result2222;
wire  [15:0] result2223;
wire  [15:0] result2224;
wire  [15:0] result2225;
wire  [15:0] result2226;
wire  [15:0] result2227;
wire  [15:0] result2228;
wire  [15:0] result2229;
wire  [15:0] result2230;
wire  [15:0] result2231;
wire  [15:0] result2232;
wire  [15:0] result2233;
wire  [15:0] result2234;
wire  [15:0] result2235;
wire  [15:0] result2236;
wire  [15:0] result2237;
wire  [15:0] result2238;
wire  [15:0] result2239;
wire  [15:0] result2240;
wire  [15:0] result2241;
wire  [15:0] result2242;
wire  [15:0] result2243;
wire  [15:0] result2244;
wire  [15:0] result2245;
wire  [15:0] result2246;
wire  [15:0] result2247;
wire  [15:0] result2248;
wire  [15:0] result2249;
wire  [15:0] result2250;
wire  [15:0] result2251;
wire  [15:0] result2252;
wire  [15:0] result2253;
wire  [15:0] result2254;
wire  [15:0] result2255;
wire  [15:0] result2256;
wire  [15:0] result2257;
wire  [15:0] result2258;
wire  [15:0] result2259;
wire  [15:0] result2260;
wire  [15:0] result2261;
wire  [15:0] result2262;
wire  [15:0] result2263;
wire  [15:0] result2264;
wire  [15:0] result2265;
wire  [15:0] result2266;
wire  [15:0] result2267;
wire  [15:0] result2268;
wire  [15:0] result2269;
wire  [15:0] result2270;
wire  [15:0] result2271;
wire  [15:0] result2272;
wire  [15:0] result2273;
wire  [15:0] result2274;
wire  [15:0] result2275;
wire  [15:0] result2276;
wire  [15:0] result2277;
wire  [15:0] result2278;
wire  [15:0] result2279;
wire  [15:0] result2280;
wire  [15:0] result2281;
wire  [15:0] result2282;
wire  [15:0] result2283;
wire  [15:0] result2284;
wire  [15:0] result2285;
wire  [15:0] result2286;
wire  [15:0] result2287;
wire  [15:0] result2288;
wire  [15:0] result2289;
wire  [15:0] result2290;
wire  [15:0] result2291;
wire  [15:0] result2292;
wire  [15:0] result2293;
wire  [15:0] result2294;
wire  [15:0] result2295;
wire  [15:0] result2296;
wire  [15:0] result2297;
wire  [15:0] result2298;
wire  [15:0] result2299;
wire  [15:0] result2300;
wire  [15:0] result2301;
wire  [15:0] result2302;
wire  [15:0] result2303;
wire  [15:0] result2304;
wire  [15:0] result2305;
wire  [15:0] result2306;
wire  [15:0] result2307;
wire  [15:0] result2308;
wire  [15:0] result2309;
wire  [15:0] result2310;
wire  [15:0] result2311;
wire  [15:0] result2312;
wire  [15:0] result2313;
wire  [15:0] result2314;
wire  [15:0] result2315;
wire  [15:0] result2316;
wire  [15:0] result2317;
wire  [15:0] result2318;
wire  [15:0] result2319;
wire  [15:0] result2320;
wire  [15:0] result2321;
wire  [15:0] result2322;
wire  [15:0] result2323;
wire  [15:0] result2324;
wire  [15:0] result2325;
wire  [15:0] result2326;
wire  [15:0] result2327;
wire  [15:0] result2328;
wire  [15:0] result2329;
wire  [15:0] result2330;
wire  [15:0] result2331;
wire  [15:0] result2332;
wire  [15:0] result2333;
wire  [15:0] result2334;
wire  [15:0] result2335;
wire  [15:0] result2336;
wire  [15:0] result2337;
wire  [15:0] result2338;
wire  [15:0] result2339;
wire  [15:0] result2340;
wire  [15:0] result2341;
wire  [15:0] result2342;
wire  [15:0] result2343;
wire  [15:0] result2344;
wire  [15:0] result2345;
wire  [15:0] result2346;
wire  [15:0] result2347;
wire  [15:0] result2348;
wire  [15:0] result2349;
wire  [15:0] result2350;
wire  [15:0] result2351;
wire  [15:0] result2352;
wire  [15:0] result2353;
wire  [15:0] result2354;
wire  [15:0] result2355;
wire  [15:0] result2356;
wire  [15:0] result2357;
wire  [15:0] result2358;
wire  [15:0] result2359;
wire  [15:0] result2360;
wire  [15:0] result2361;
wire  [15:0] result2362;
wire  [15:0] result2363;
wire  [15:0] result2364;
wire  [15:0] result2365;
wire  [15:0] result2366;
wire  [15:0] result2367;
wire  [15:0] result2368;
wire  [15:0] result2369;
wire  [15:0] result2370;
wire  [15:0] result2371;
wire  [15:0] result2372;
wire  [15:0] result2373;
wire  [15:0] result2374;
wire  [15:0] result2375;
wire  [15:0] result2376;
wire  [15:0] result2377;
wire  [15:0] result2378;
wire  [15:0] result2379;
wire  [15:0] result2380;
wire  [15:0] result2381;
wire  [15:0] result2382;
wire  [15:0] result2383;
wire  [15:0] result2384;
wire  [15:0] result2385;
wire  [15:0] result2386;
wire  [15:0] result2387;
wire  [15:0] result2388;
wire  [15:0] result2389;
wire  [15:0] result2390;
wire  [15:0] result2391;
wire  [15:0] result2392;
wire  [15:0] result2393;
wire  [15:0] result2394;
wire  [15:0] result2395;
wire  [15:0] result2396;
wire  [15:0] result2397;
wire  [15:0] result2398;
wire  [15:0] result2399;
wire  [15:0] result2400;
wire  [15:0] result2401;
wire  [15:0] result2402;
wire  [15:0] result2403;
wire  [15:0] result2404;
wire  [15:0] result2405;
wire  [15:0] result2406;
wire  [15:0] result2407;
wire  [15:0] result2408;
wire  [15:0] result2409;
wire  [15:0] result2410;
wire  [15:0] result2411;
wire  [15:0] result2412;
wire  [15:0] result2413;
wire  [15:0] result2414;
wire  [15:0] result2415;
wire  [15:0] result2416;
wire  [15:0] result2417;
wire  [15:0] result2418;
wire  [15:0] result2419;
wire  [15:0] result2420;
wire  [15:0] result2421;
wire  [15:0] result2422;
wire  [15:0] result2423;
wire  [15:0] result2424;
wire  [15:0] result2425;
wire  [15:0] result2426;
wire  [15:0] result2427;
wire  [15:0] result2428;
wire  [15:0] result2429;
wire  [15:0] result2430;
wire  [15:0] result2431;
wire  [15:0] result2432;
wire  [15:0] result2433;
wire  [15:0] result2434;
wire  [15:0] result2435;
wire  [15:0] result2436;
wire  [15:0] result2437;
wire  [15:0] result2438;
wire  [15:0] result2439;
wire  [15:0] result2440;
wire  [15:0] result2441;
wire  [15:0] result2442;
wire  [15:0] result2443;
wire  [15:0] result2444;
wire  [15:0] result2445;
wire  [15:0] result2446;
wire  [15:0] result2447;
wire  [15:0] result2448;
wire  [15:0] result2449;
wire  [15:0] result2450;
wire  [15:0] result2451;
wire  [15:0] result2452;
wire  [15:0] result2453;
wire  [15:0] result2454;
wire  [15:0] result2455;
wire  [15:0] result2456;
wire  [15:0] result2457;
wire  [15:0] result2458;
wire  [15:0] result2459;
wire  [15:0] result2460;
wire  [15:0] result2461;
wire  [15:0] result2462;
wire  [15:0] result2463;
wire  [15:0] result2464;
wire  [15:0] result2465;
wire  [15:0] result2466;
wire  [15:0] result2467;
wire  [15:0] result2468;
wire  [15:0] result2469;
wire  [15:0] result2470;
wire  [15:0] result2471;
wire  [15:0] result2472;
wire  [15:0] result2473;
wire  [15:0] result2474;
wire  [15:0] result2475;
wire  [15:0] result2476;
wire  [15:0] result2477;
wire  [15:0] result2478;
wire  [15:0] result2479;
wire  [15:0] result2480;
wire  [15:0] result2481;
wire  [15:0] result2482;
wire  [15:0] result2483;
wire  [15:0] result2484;
wire  [15:0] result2485;
wire  [15:0] result2486;
wire  [15:0] result2487;
wire  [15:0] result2488;
wire  [15:0] result2489;
wire  [15:0] result2490;
wire  [15:0] result2491;
wire  [15:0] result2492;
wire  [15:0] result2493;
wire  [15:0] result2494;
wire  [15:0] result2495;
wire  [15:0] result2496;
wire  [15:0] result2497;
wire  [15:0] result2498;
wire  [15:0] result2499;
wire  [15:0] result2500;
wire  [15:0] result2501;
wire  [15:0] result2502;
wire  [15:0] result2503;
wire  [15:0] result2504;
wire  [15:0] result2505;
wire  [15:0] result2506;
wire  [15:0] result2507;
wire  [15:0] result2508;
wire  [15:0] result2509;
wire  [15:0] result2510;
wire  [15:0] result2511;
wire  [15:0] result2512;
wire  [15:0] result2513;
wire  [15:0] result2514;
wire  [15:0] result2515;
wire  [15:0] result2516;
wire  [15:0] result2517;
wire  [15:0] result2518;
wire  [15:0] result2519;
wire  [15:0] result2520;
wire  [15:0] result2521;
wire  [15:0] result2522;
wire  [15:0] result2523;
wire  [15:0] result2524;
wire  [15:0] result2525;
wire  [15:0] result2526;
wire  [15:0] result2527;
wire  [15:0] result2528;
wire  [15:0] result2529;
wire  [15:0] result2530;
wire  [15:0] result2531;
wire  [15:0] result2532;
wire  [15:0] result2533;
wire  [15:0] result2534;
wire  [15:0] result2535;
wire  [15:0] result2536;
wire  [15:0] result2537;
wire  [15:0] result2538;
wire  [15:0] result2539;
wire  [15:0] result2540;
wire  [15:0] result2541;
wire  [15:0] result2542;
wire  [15:0] result2543;
wire  [15:0] result2544;
wire  [15:0] result2545;
wire  [15:0] result2546;
wire  [15:0] result2547;
wire  [15:0] result2548;
wire  [15:0] result2549;
wire  [15:0] result2550;
wire  [15:0] result2551;
wire  [15:0] result2552;
wire  [15:0] result2553;
wire  [15:0] result2554;
wire  [15:0] result2555;
wire  [15:0] result2556;
wire  [15:0] result2557;
wire  [15:0] result2558;
wire  [15:0] result2559;
wire  [15:0] result2560;
wire  [15:0] result2561;
wire  [15:0] result2562;
wire  [15:0] result2563;
wire  [15:0] result2564;
wire  [15:0] result2565;
wire  [15:0] result2566;
wire  [15:0] result2567;
wire  [15:0] result2568;
wire  [15:0] result2569;
wire  [15:0] result2570;
wire  [15:0] result2571;
wire  [15:0] result2572;
wire  [15:0] result2573;
wire  [15:0] result2574;
wire  [15:0] result2575;
wire  [15:0] result2576;
wire  [15:0] result2577;
wire  [15:0] result2578;
wire  [15:0] result2579;
wire  [15:0] result2580;
wire  [15:0] result2581;
wire  [15:0] result2582;
wire  [15:0] result2583;
wire  [15:0] result2584;
wire  [15:0] result2585;
wire  [15:0] result2586;
wire  [15:0] result2587;
wire  [15:0] result2588;
wire  [15:0] result2589;
wire  [15:0] result2590;
wire  [15:0] result2591;
wire  [15:0] result2592;
wire  [15:0] result2593;
wire  [15:0] result2594;
wire  [15:0] result2595;
wire  [15:0] result2596;
wire  [15:0] result2597;
wire  [15:0] result2598;
wire  [15:0] result2599;
wire  [15:0] result2600;
wire  [15:0] result2601;
wire  [15:0] result2602;
wire  [15:0] result2603;
wire  [15:0] result2604;
wire  [15:0] result2605;
wire  [15:0] result2606;
wire  [15:0] result2607;
wire  [15:0] result2608;
wire  [15:0] result2609;
wire  [15:0] result2610;
wire  [15:0] result2611;
wire  [15:0] result2612;
wire  [15:0] result2613;
wire  [15:0] result2614;
wire  [15:0] result2615;
wire  [15:0] result2616;
wire  [15:0] result2617;
wire  [15:0] result2618;
wire  [15:0] result2619;
wire  [15:0] result2620;
wire  [15:0] result2621;
wire  [15:0] result2622;
wire  [15:0] result2623;
wire  [15:0] result2624;
wire  [15:0] result2625;
wire  [15:0] result2626;
wire  [15:0] result2627;
wire  [15:0] result2628;
wire  [15:0] result2629;
wire  [15:0] result2630;
wire  [15:0] result2631;
wire  [15:0] result2632;
wire  [15:0] result2633;
wire  [15:0] result2634;
wire  [15:0] result2635;
wire  [15:0] result2636;
wire  [15:0] result2637;
wire  [15:0] result2638;
wire  [15:0] result2639;
wire  [15:0] result2640;
wire  [15:0] result2641;
wire  [15:0] result2642;
wire  [15:0] result2643;
wire  [15:0] result2644;
wire  [15:0] result2645;
wire  [15:0] result2646;
wire  [15:0] result2647;
wire  [15:0] result2648;
wire  [15:0] result2649;
wire  [15:0] result2650;
wire  [15:0] result2651;
wire  [15:0] result2652;
wire  [15:0] result2653;
wire  [15:0] result2654;
wire  [15:0] result2655;
wire  [15:0] result2656;
wire  [15:0] result2657;
wire  [15:0] result2658;
wire  [15:0] result2659;
wire  [15:0] result2660;
wire  [15:0] result2661;
wire  [15:0] result2662;
wire  [15:0] result2663;
wire  [15:0] result2664;
wire  [15:0] result2665;
wire  [15:0] result2666;
wire  [15:0] result2667;
wire  [15:0] result2668;
wire  [15:0] result2669;
wire  [15:0] result2670;
wire  [15:0] result2671;
wire  [15:0] result2672;
wire  [15:0] result2673;
wire  [15:0] result2674;
wire  [15:0] result2675;
wire  [15:0] result2676;
wire  [15:0] result2677;
wire  [15:0] result2678;
wire  [15:0] result2679;
wire  [15:0] result2680;
wire  [15:0] result2681;
wire  [15:0] result2682;
wire  [15:0] result2683;
wire  [15:0] result2684;
wire  [15:0] result2685;
wire  [15:0] result2686;
wire  [15:0] result2687;
wire  [15:0] result2688;
wire  [15:0] result2689;
wire  [15:0] result2690;
wire  [15:0] result2691;
wire  [15:0] result2692;
wire  [15:0] result2693;
wire  [15:0] result2694;
wire  [15:0] result2695;
wire  [15:0] result2696;
wire  [15:0] result2697;
wire  [15:0] result2698;
wire  [15:0] result2699;
wire  [15:0] result2700;
wire  [15:0] result2701;
wire  [15:0] result2702;
wire  [15:0] result2703;
wire  [15:0] result2704;
wire  [15:0] result2705;
wire  [15:0] result2706;
wire  [15:0] result2707;
wire  [15:0] result2708;
wire  [15:0] result2709;
wire  [15:0] result2710;
wire  [15:0] result2711;
wire  [15:0] result2712;
wire  [15:0] result2713;
wire  [15:0] result2714;
wire  [15:0] result2715;
wire  [15:0] result2716;
wire  [15:0] result2717;
wire  [15:0] result2718;
wire  [15:0] result2719;
wire  [15:0] result2720;
wire  [15:0] result2721;
wire  [15:0] result2722;
wire  [15:0] result2723;
wire  [15:0] result2724;
wire  [15:0] result2725;
wire  [15:0] result2726;
wire  [15:0] result2727;
wire  [15:0] result2728;
wire  [15:0] result2729;
wire  [15:0] result2730;
wire  [15:0] result2731;
wire  [15:0] result2732;
wire  [15:0] result2733;
wire  [15:0] result2734;
wire  [15:0] result2735;
wire  [15:0] result2736;
wire  [15:0] result2737;
wire  [15:0] result2738;
wire  [15:0] result2739;
wire  [15:0] result2740;
wire  [15:0] result2741;
wire  [15:0] result2742;
wire  [15:0] result2743;
wire  [15:0] result2744;
wire  [15:0] result2745;
wire  [15:0] result2746;
wire  [15:0] result2747;
wire  [15:0] result2748;
wire  [15:0] result2749;
wire  [15:0] result2750;
wire  [15:0] result2751;
wire  [15:0] result2752;
wire  [15:0] result2753;
wire  [15:0] result2754;
wire  [15:0] result2755;
wire  [15:0] result2756;
wire  [15:0] result2757;
wire  [15:0] result2758;
wire  [15:0] result2759;
wire  [15:0] result2760;
wire  [15:0] result2761;
wire  [15:0] result2762;
wire  [15:0] result2763;
wire  [15:0] result2764;
wire  [15:0] result2765;
wire  [15:0] result2766;
wire  [15:0] result2767;
wire  [15:0] result2768;
wire  [15:0] result2769;
wire  [15:0] result2770;
wire  [15:0] result2771;
wire  [15:0] result2772;
wire  [15:0] result2773;
wire  [15:0] result2774;
wire  [15:0] result2775;
wire  [15:0] result2776;
wire  [15:0] result2777;
wire  [15:0] result2778;
wire  [15:0] result2779;
wire  [15:0] result2780;
wire  [15:0] result2781;
wire  [15:0] result2782;
wire  [15:0] result2783;
wire  [15:0] result2784;
wire  [15:0] result2785;
wire  [15:0] result2786;
wire  [15:0] result2787;
wire  [15:0] result2788;
wire  [15:0] result2789;
wire  [15:0] result2790;
wire  [15:0] result2791;
wire  [15:0] result2792;
wire  [15:0] result2793;
wire  [15:0] result2794;
wire  [15:0] result2795;
wire  [15:0] result2796;
wire  [15:0] result2797;
wire  [15:0] result2798;
wire  [15:0] result2799;
wire  [15:0] result2800;
wire  [15:0] result2801;
wire  [15:0] result2802;
wire  [15:0] result2803;
wire  [15:0] result2804;
wire  [15:0] result2805;
wire  [15:0] result2806;
wire  [15:0] result2807;
wire  [15:0] result2808;
wire  [15:0] result2809;
wire  [15:0] result2810;
wire  [15:0] result2811;
wire  [15:0] result2812;
wire  [15:0] result2813;
wire  [15:0] result2814;
wire  [15:0] result2815;
wire  [15:0] result2816;
wire  [15:0] result2817;
wire  [15:0] result2818;
wire  [15:0] result2819;
wire  [15:0] result2820;
wire  [15:0] result2821;
wire  [15:0] result2822;
wire  [15:0] result2823;
wire  [15:0] result2824;
wire  [15:0] result2825;
wire  [15:0] result2826;
wire  [15:0] result2827;
wire  [15:0] result2828;
wire  [15:0] result2829;
wire  [15:0] result2830;
wire  [15:0] result2831;
wire  [15:0] result2832;
wire  [15:0] result2833;
wire  [15:0] result2834;
wire  [15:0] result2835;
wire  [15:0] result2836;
wire  [15:0] result2837;
wire  [15:0] result2838;
wire  [15:0] result2839;
wire  [15:0] result2840;
wire  [15:0] result2841;
wire  [15:0] result2842;
wire  [15:0] result2843;
wire  [15:0] result2844;
wire  [15:0] result2845;
wire  [15:0] result2846;
wire  [15:0] result2847;
wire  [15:0] result2848;
wire  [15:0] result2849;
wire  [15:0] result2850;
wire  [15:0] result2851;
wire  [15:0] result2852;
wire  [15:0] result2853;
wire  [15:0] result2854;
wire  [15:0] result2855;
wire  [15:0] result2856;
wire  [15:0] result2857;
wire  [15:0] result2858;
wire  [15:0] result2859;
wire  [15:0] result2860;
wire  [15:0] result2861;
wire  [15:0] result2862;
wire  [15:0] result2863;
wire  [15:0] result2864;
wire  [15:0] result2865;
wire  [15:0] result2866;
wire  [15:0] result2867;
wire  [15:0] result2868;
wire  [15:0] result2869;
wire  [15:0] result2870;
wire  [15:0] result2871;
wire  [15:0] result2872;
wire  [15:0] result2873;
wire  [15:0] result2874;
wire  [15:0] result2875;
wire  [15:0] result2876;
wire  [15:0] result2877;
wire  [15:0] result2878;
wire  [15:0] result2879;
wire  [15:0] result2880;
wire  [15:0] result2881;
wire  [15:0] result2882;
wire  [15:0] result2883;
wire  [15:0] result2884;
wire  [15:0] result2885;
wire  [15:0] result2886;
wire  [15:0] result2887;
wire  [15:0] result2888;
wire  [15:0] result2889;
wire  [15:0] result2890;
wire  [15:0] result2891;
wire  [15:0] result2892;
wire  [15:0] result2893;
wire  [15:0] result2894;
wire  [15:0] result2895;
wire  [15:0] result2896;
wire  [15:0] result2897;
wire  [15:0] result2898;
wire  [15:0] result2899;
wire  [15:0] result2900;
wire  [15:0] result2901;
wire  [15:0] result2902;
wire  [15:0] result2903;
wire  [15:0] result2904;
wire  [15:0] result2905;
wire  [15:0] result2906;
wire  [15:0] result2907;
wire  [15:0] result2908;
wire  [15:0] result2909;
wire  [15:0] result2910;
wire  [15:0] result2911;
wire  [15:0] result2912;
wire  [15:0] result2913;
wire  [15:0] result2914;
wire  [15:0] result2915;
wire  [15:0] result2916;
wire  [15:0] result2917;
wire  [15:0] result2918;
wire  [15:0] result2919;
wire  [15:0] result2920;
wire  [15:0] result2921;
wire  [15:0] result2922;
wire  [15:0] result2923;
wire  [15:0] result2924;
wire  [15:0] result2925;
wire  [15:0] result2926;
wire  [15:0] result2927;
wire  [15:0] result2928;
wire  [15:0] result2929;
wire  [15:0] result2930;
wire  [15:0] result2931;
wire  [15:0] result2932;
wire  [15:0] result2933;
wire  [15:0] result2934;
wire  [15:0] result2935;
wire  [15:0] result2936;
wire  [15:0] result2937;
wire  [15:0] result2938;
wire  [15:0] result2939;
wire  [15:0] result2940;
wire  [15:0] result2941;
wire  [15:0] result2942;
wire  [15:0] result2943;
wire  [15:0] result2944;
wire  [15:0] result2945;
wire  [15:0] result2946;
wire  [15:0] result2947;
wire  [15:0] result2948;
wire  [15:0] result2949;
wire  [15:0] result2950;
wire  [15:0] result2951;
wire  [15:0] result2952;
wire  [15:0] result2953;
wire  [15:0] result2954;
wire  [15:0] result2955;
wire  [15:0] result2956;
wire  [15:0] result2957;
wire  [15:0] result2958;
wire  [15:0] result2959;
wire  [15:0] result2960;
wire  [15:0] result2961;
wire  [15:0] result2962;
wire  [15:0] result2963;
wire  [15:0] result2964;
wire  [15:0] result2965;
wire  [15:0] result2966;
wire  [15:0] result2967;
wire  [15:0] result2968;
wire  [15:0] result2969;
wire  [15:0] result2970;
wire  [15:0] result2971;
wire  [15:0] result2972;
wire  [15:0] result2973;
wire  [15:0] result2974;
wire  [15:0] result2975;
wire  [15:0] result2976;
wire  [15:0] result2977;
wire  [15:0] result2978;
wire  [15:0] result2979;
wire  [15:0] result2980;
wire  [15:0] result2981;
wire  [15:0] result2982;
wire  [15:0] result2983;
wire  [15:0] result2984;
wire  [15:0] result2985;
wire  [15:0] result2986;
wire  [15:0] result2987;
wire  [15:0] result2988;
wire  [15:0] result2989;
wire  [15:0] result2990;
wire  [15:0] result2991;
wire  [15:0] result2992;
wire  [15:0] result2993;
wire  [15:0] result2994;
wire  [15:0] result2995;
wire  [15:0] result2996;
wire  [15:0] result2997;
wire  [15:0] result2998;
wire  [15:0] result2999;
wire  [15:0] result3000;
wire  [15:0] result3001;
wire  [15:0] result3002;
wire  [15:0] result3003;
wire  [15:0] result3004;
wire  [15:0] result3005;
wire  [15:0] result3006;
wire  [15:0] result3007;
wire  [15:0] result3008;
wire  [15:0] result3009;
wire  [15:0] result3010;
wire  [15:0] result3011;
wire  [15:0] result3012;
wire  [15:0] result3013;
wire  [15:0] result3014;
wire  [15:0] result3015;
wire  [15:0] result3016;
wire  [15:0] result3017;
wire  [15:0] result3018;
wire  [15:0] result3019;
wire  [15:0] result3020;
wire  [15:0] result3021;
wire  [15:0] result3022;
wire  [15:0] result3023;
wire  [15:0] result3024;
wire  [15:0] result3025;
wire  [15:0] result3026;
wire  [15:0] result3027;
wire  [15:0] result3028;
wire  [15:0] result3029;
wire  [15:0] result3030;
wire  [15:0] result3031;
wire  [15:0] result3032;
wire  [15:0] result3033;
wire  [15:0] result3034;
wire  [15:0] result3035;
wire  [15:0] result3036;
wire  [15:0] result3037;
wire  [15:0] result3038;
wire  [15:0] result3039;
wire  [15:0] result3040;
wire  [15:0] result3041;
wire  [15:0] result3042;
wire  [15:0] result3043;
wire  [15:0] result3044;
wire  [15:0] result3045;
wire  [15:0] result3046;
wire  [15:0] result3047;
wire  [15:0] result3048;
wire  [15:0] result3049;
wire  [15:0] result3050;
wire  [15:0] result3051;
wire  [15:0] result3052;
wire  [15:0] result3053;
wire  [15:0] result3054;
wire  [15:0] result3055;
wire  [15:0] result3056;
wire  [15:0] result3057;
wire  [15:0] result3058;
wire  [15:0] result3059;
wire  [15:0] result3060;
wire  [15:0] result3061;
wire  [15:0] result3062;
wire  [15:0] result3063;
wire  [15:0] result3064;
wire  [15:0] result3065;
wire  [15:0] result3066;
wire  [15:0] result3067;
wire  [15:0] result3068;
wire  [15:0] result3069;
wire  [15:0] result3070;
wire  [15:0] result3071;
wire  [15:0] result3072;
wire  [15:0] result3073;
wire  [15:0] result3074;
wire  [15:0] result3075;
wire  [15:0] result3076;
wire  [15:0] result3077;
wire  [15:0] result3078;
wire  [15:0] result3079;
wire  [15:0] result3080;
wire  [15:0] result3081;
wire  [15:0] result3082;
wire  [15:0] result3083;
wire  [15:0] result3084;
wire  [15:0] result3085;
wire  [15:0] result3086;
wire  [15:0] result3087;
wire  [15:0] result3088;
wire  [15:0] result3089;
wire  [15:0] result3090;
wire  [15:0] result3091;
wire  [15:0] result3092;
wire  [15:0] result3093;
wire  [15:0] result3094;
wire  [15:0] result3095;
wire  [15:0] result3096;
wire  [15:0] result3097;
wire  [15:0] result3098;
wire  [15:0] result3099;
wire  [15:0] result3100;
wire  [15:0] result3101;
wire  [15:0] result3102;
wire  [15:0] result3103;
wire  [15:0] result3104;
wire  [15:0] result3105;
wire  [15:0] result3106;
wire  [15:0] result3107;
wire  [15:0] result3108;
wire  [15:0] result3109;
wire  [15:0] result3110;
wire  [15:0] result3111;
wire  [15:0] result3112;
wire  [15:0] result3113;
wire  [15:0] result3114;
wire  [15:0] result3115;
wire  [15:0] result3116;
wire  [15:0] result3117;
wire  [15:0] result3118;
wire  [15:0] result3119;
wire  [15:0] result3120;
wire  [15:0] result3121;
wire  [15:0] result3122;
wire  [15:0] result3123;
wire  [15:0] result3124;
wire  [15:0] result3125;
wire  [15:0] result3126;
wire  [15:0] result3127;
wire  [15:0] result3128;
wire  [15:0] result3129;
wire  [15:0] result3130;
wire  [15:0] result3131;
wire  [15:0] result3132;
wire  [15:0] result3133;
wire  [15:0] result3134;
wire  [15:0] result3135;
wire  [15:0] result3136;
wire  [15:0] result3137;
wire  [15:0] result3138;
wire  [15:0] result3139;
wire  [15:0] result3140;
wire  [15:0] result3141;
wire  [15:0] result3142;
wire  [15:0] result3143;
wire  [15:0] result3144;
wire  [15:0] result3145;
wire  [15:0] result3146;
wire  [15:0] result3147;
wire  [15:0] result3148;
wire  [15:0] result3149;
wire  [15:0] result3150;
wire  [15:0] result3151;
wire  [15:0] result3152;
wire  [15:0] result3153;
wire  [15:0] result3154;
wire  [15:0] result3155;
wire  [15:0] result3156;
wire  [15:0] result3157;
wire  [15:0] result3158;
wire  [15:0] result3159;
wire  [15:0] result3160;
wire  [15:0] result3161;
wire  [15:0] result3162;
wire  [15:0] result3163;
wire  [15:0] result3164;
wire  [15:0] result3165;
wire  [15:0] result3166;
wire  [15:0] result3167;
wire  [15:0] result3168;
wire  [15:0] result3169;
wire  [15:0] result3170;
wire  [15:0] result3171;
wire  [15:0] result3172;
wire  [15:0] result3173;
wire  [15:0] result3174;
wire  [15:0] result3175;
wire  [15:0] result3176;
wire  [15:0] result3177;
wire  [15:0] result3178;
wire  [15:0] result3179;
wire  [15:0] result3180;
wire  [15:0] result3181;
wire  [15:0] result3182;
wire  [15:0] result3183;
wire  [15:0] result3184;
wire  [15:0] result3185;
wire  [15:0] result3186;
wire  [15:0] result3187;
wire  [15:0] result3188;
wire  [15:0] result3189;
wire  [15:0] result3190;
wire  [15:0] result3191;
wire  [15:0] result3192;
wire  [15:0] result3193;
wire  [15:0] result3194;
wire  [15:0] result3195;
wire  [15:0] result3196;
wire  [15:0] result3197;
wire  [15:0] result3198;
wire  [15:0] result3199;
wire  [15:0] result3200;
wire  [15:0] result3201;
wire  [15:0] result3202;
wire  [15:0] result3203;
wire  [15:0] result3204;
wire  [15:0] result3205;
wire  [15:0] result3206;
wire  [15:0] result3207;
wire  [15:0] result3208;
wire  [15:0] result3209;
wire  [15:0] result3210;
wire  [15:0] result3211;
wire  [15:0] result3212;
wire  [15:0] result3213;
wire  [15:0] result3214;
wire  [15:0] result3215;
wire  [15:0] result3216;
wire  [15:0] result3217;
wire  [15:0] result3218;
wire  [15:0] result3219;
wire  [15:0] result3220;
wire  [15:0] result3221;
wire  [15:0] result3222;
wire  [15:0] result3223;
wire  [15:0] result3224;
wire  [15:0] result3225;
wire  [15:0] result3226;
wire  [15:0] result3227;
wire  [15:0] result3228;
wire  [15:0] result3229;
wire  [15:0] result3230;
wire  [15:0] result3231;
wire  [15:0] result3232;
wire  [15:0] result3233;
wire  [15:0] result3234;
wire  [15:0] result3235;
wire  [15:0] result3236;
wire  [15:0] result3237;
wire  [15:0] result3238;
wire  [15:0] result3239;
wire  [15:0] result3240;
wire  [15:0] result3241;
wire  [15:0] result3242;
wire  [15:0] result3243;
wire  [15:0] result3244;
wire  [15:0] result3245;
wire  [15:0] result3246;
wire  [15:0] result3247;
wire  [15:0] result3248;
wire  [15:0] result3249;
wire  [15:0] result3250;
wire  [15:0] result3251;
wire  [15:0] result3252;
wire  [15:0] result3253;
wire  [15:0] result3254;
wire  [15:0] result3255;
wire  [15:0] result3256;
wire  [15:0] result3257;
wire  [15:0] result3258;
wire  [15:0] result3259;
wire  [15:0] result3260;
wire  [15:0] result3261;
wire  [15:0] result3262;
wire  [15:0] result3263;
wire  [15:0] result3264;
wire  [15:0] result3265;
wire  [15:0] result3266;
wire  [15:0] result3267;
wire  [15:0] result3268;
wire  [15:0] result3269;
wire  [15:0] result3270;
wire  [15:0] result3271;
wire  [15:0] result3272;
wire  [15:0] result3273;
wire  [15:0] result3274;
wire  [15:0] result3275;
wire  [15:0] result3276;
wire  [15:0] result3277;
wire  [15:0] result3278;
wire  [15:0] result3279;
wire  [15:0] result3280;
wire  [15:0] result3281;
wire  [15:0] result3282;
wire  [15:0] result3283;
wire  [15:0] result3284;
wire  [15:0] result3285;
wire  [15:0] result3286;
wire  [15:0] result3287;
wire  [15:0] result3288;
wire  [15:0] result3289;
wire  [15:0] result3290;
wire  [15:0] result3291;
wire  [15:0] result3292;
wire  [15:0] result3293;
wire  [15:0] result3294;
wire  [15:0] result3295;
wire  [15:0] result3296;
wire  [15:0] result3297;
wire  [15:0] result3298;
wire  [15:0] result3299;
wire  [15:0] result3300;
wire  [15:0] result3301;
wire  [15:0] result3302;
wire  [15:0] result3303;
wire  [15:0] result3304;
wire  [15:0] result3305;
wire  [15:0] result3306;
wire  [15:0] result3307;
wire  [15:0] result3308;
wire  [15:0] result3309;
wire  [15:0] result3310;
wire  [15:0] result3311;
wire  [15:0] result3312;
wire  [15:0] result3313;
wire  [15:0] result3314;
wire  [15:0] result3315;
wire  [15:0] result3316;
wire  [15:0] result3317;
wire  [15:0] result3318;
wire  [15:0] result3319;
wire  [15:0] result3320;
wire  [15:0] result3321;
wire  [15:0] result3322;
wire  [15:0] result3323;
wire  [15:0] result3324;
wire  [15:0] result3325;
wire  [15:0] result3326;
wire  [15:0] result3327;
wire  [15:0] result3328;
wire  [15:0] result3329;
wire  [15:0] result3330;
wire  [15:0] result3331;
wire  [15:0] result3332;
wire  [15:0] result3333;
wire  [15:0] result3334;
wire  [15:0] result3335;
wire  [15:0] result3336;
wire  [15:0] result3337;
wire  [15:0] result3338;
wire  [15:0] result3339;
wire  [15:0] result3340;
wire  [15:0] result3341;
wire  [15:0] result3342;
wire  [15:0] result3343;
wire  [15:0] result3344;
wire  [15:0] result3345;
wire  [15:0] result3346;
wire  [15:0] result3347;
wire  [15:0] result3348;
wire  [15:0] result3349;
wire  [15:0] result3350;
wire  [15:0] result3351;
wire  [15:0] result3352;
wire  [15:0] result3353;
wire  [15:0] result3354;
wire  [15:0] result3355;
wire  [15:0] result3356;
wire  [15:0] result3357;
wire  [15:0] result3358;
wire  [15:0] result3359;
wire  [15:0] result3360;
wire  [15:0] result3361;
wire  [15:0] result3362;
wire  [15:0] result3363;
wire  [15:0] result3364;
wire  [15:0] result3365;
wire  [15:0] result3366;
wire  [15:0] result3367;
wire  [15:0] result3368;
wire  [15:0] result3369;
wire  [15:0] result3370;
wire  [15:0] result3371;
wire  [15:0] result3372;
wire  [15:0] result3373;
wire  [15:0] result3374;
wire  [15:0] result3375;
wire  [15:0] result3376;
wire  [15:0] result3377;
wire  [15:0] result3378;
wire  [15:0] result3379;
wire  [15:0] result3380;
wire  [15:0] result3381;
wire  [15:0] result3382;
wire  [15:0] result3383;
wire  [15:0] result3384;
wire  [15:0] result3385;
wire  [15:0] result3386;
wire  [15:0] result3387;
wire  [15:0] result3388;
wire  [15:0] result3389;
wire  [15:0] result3390;
wire  [15:0] result3391;
wire  [15:0] result3392;
wire  [15:0] result3393;
wire  [15:0] result3394;
wire  [15:0] result3395;
wire  [15:0] result3396;
wire  [15:0] result3397;
wire  [15:0] result3398;
wire  [15:0] result3399;
wire  [15:0] result3400;
wire  [15:0] result3401;
wire  [15:0] result3402;
wire  [15:0] result3403;
wire  [15:0] result3404;
wire  [15:0] result3405;
wire  [15:0] result3406;
wire  [15:0] result3407;
wire  [15:0] result3408;
wire  [15:0] result3409;
wire  [15:0] result3410;
wire  [15:0] result3411;
wire  [15:0] result3412;
wire  [15:0] result3413;
wire  [15:0] result3414;
wire  [15:0] result3415;
wire  [15:0] result3416;
wire  [15:0] result3417;
wire  [15:0] result3418;
wire  [15:0] result3419;
wire  [15:0] result3420;
wire  [15:0] result3421;
wire  [15:0] result3422;
wire  [15:0] result3423;
wire  [15:0] result3424;
wire  [15:0] result3425;
wire  [15:0] result3426;
wire  [15:0] result3427;
wire  [15:0] result3428;
wire  [15:0] result3429;
wire  [15:0] result3430;
wire  [15:0] result3431;
wire  [15:0] result3432;
wire  [15:0] result3433;
wire  [15:0] result3434;
wire  [15:0] result3435;
wire  [15:0] result3436;
wire  [15:0] result3437;
wire  [15:0] result3438;
wire  [15:0] result3439;
wire  [15:0] result3440;
wire  [15:0] result3441;
wire  [15:0] result3442;
wire  [15:0] result3443;
wire  [15:0] result3444;
wire  [15:0] result3445;
wire  [15:0] result3446;
wire  [15:0] result3447;
wire  [15:0] result3448;
wire  [15:0] result3449;
wire  [15:0] result3450;
wire  [15:0] result3451;
wire  [15:0] result3452;
wire  [15:0] result3453;
wire  [15:0] result3454;
wire  [15:0] result3455;
wire  [15:0] result3456;
wire  [15:0] result3457;
wire  [15:0] result3458;
wire  [15:0] result3459;
wire  [15:0] result3460;
wire  [15:0] result3461;
wire  [15:0] result3462;
wire  [15:0] result3463;
wire  [15:0] result3464;
wire  [15:0] result3465;
wire  [15:0] result3466;
wire  [15:0] result3467;
wire  [15:0] result3468;
wire  [15:0] result3469;
wire  [15:0] result3470;
wire  [15:0] result3471;
wire  [15:0] result3472;
wire  [15:0] result3473;
wire  [15:0] result3474;
wire  [15:0] result3475;
wire  [15:0] result3476;
wire  [15:0] result3477;
wire  [15:0] result3478;
wire  [15:0] result3479;
wire  [15:0] result3480;
wire  [15:0] result3481;
wire  [15:0] result3482;
wire  [15:0] result3483;
wire  [15:0] result3484;
wire  [15:0] result3485;
wire  [15:0] result3486;
wire  [15:0] result3487;
wire  [15:0] result3488;
wire  [15:0] result3489;
wire  [15:0] result3490;
wire  [15:0] result3491;
wire  [15:0] result3492;
wire  [15:0] result3493;
wire  [15:0] result3494;
wire  [15:0] result3495;
wire  [15:0] result3496;
wire  [15:0] result3497;
wire  [15:0] result3498;
wire  [15:0] result3499;
wire  [15:0] result3500;
wire  [15:0] result3501;
wire  [15:0] result3502;
wire  [15:0] result3503;
wire  [15:0] result3504;
wire  [15:0] result3505;
wire  [15:0] result3506;
wire  [15:0] result3507;
wire  [15:0] result3508;
wire  [15:0] result3509;
wire  [15:0] result3510;
wire  [15:0] result3511;
wire  [15:0] result3512;
wire  [15:0] result3513;
wire  [15:0] result3514;
wire  [15:0] result3515;
wire  [15:0] result3516;
wire  [15:0] result3517;
wire  [15:0] result3518;
wire  [15:0] result3519;
wire  [15:0] result3520;
wire  [15:0] result3521;
wire  [15:0] result3522;
wire  [15:0] result3523;
wire  [15:0] result3524;
wire  [15:0] result3525;
wire  [15:0] result3526;
wire  [15:0] result3527;
wire  [15:0] result3528;
wire  [15:0] result3529;
wire  [15:0] result3530;
wire  [15:0] result3531;
wire  [15:0] result3532;
wire  [15:0] result3533;
wire  [15:0] result3534;
wire  [15:0] result3535;
wire  [15:0] result3536;
wire  [15:0] result3537;
wire  [15:0] result3538;
wire  [15:0] result3539;
wire  [15:0] result3540;
wire  [15:0] result3541;
wire  [15:0] result3542;
wire  [15:0] result3543;
wire  [15:0] result3544;
wire  [15:0] result3545;
wire  [15:0] result3546;
wire  [15:0] result3547;
wire  [15:0] result3548;
wire  [15:0] result3549;
wire  [15:0] result3550;
wire  [15:0] result3551;
wire  [15:0] result3552;
wire  [15:0] result3553;
wire  [15:0] result3554;
wire  [15:0] result3555;
wire  [15:0] result3556;
wire  [15:0] result3557;
wire  [15:0] result3558;
wire  [15:0] result3559;
wire  [15:0] result3560;
wire  [15:0] result3561;
wire  [15:0] result3562;
wire  [15:0] result3563;
wire  [15:0] result3564;
wire  [15:0] result3565;
wire  [15:0] result3566;
wire  [15:0] result3567;
wire  [15:0] result3568;
wire  [15:0] result3569;
wire  [15:0] result3570;
wire  [15:0] result3571;
wire  [15:0] result3572;
wire  [15:0] result3573;
wire  [15:0] result3574;
wire  [15:0] result3575;
wire  [15:0] result3576;
wire  [15:0] result3577;
wire  [15:0] result3578;
wire  [15:0] result3579;
wire  [15:0] result3580;
wire  [15:0] result3581;
wire  [15:0] result3582;
wire  [15:0] result3583;
wire  [15:0] result3584;
wire  [15:0] result3585;
wire  [15:0] result3586;
wire  [15:0] result3587;
wire  [15:0] result3588;
wire  [15:0] result3589;
wire  [15:0] result3590;
wire  [15:0] result3591;
wire  [15:0] result3592;
wire  [15:0] result3593;
wire  [15:0] result3594;
wire  [15:0] result3595;
wire  [15:0] result3596;
wire  [15:0] result3597;
wire  [15:0] result3598;
wire  [15:0] result3599;
wire  [15:0] result3600;
wire  [15:0] result3601;
wire  [15:0] result3602;
wire  [15:0] result3603;
wire  [15:0] result3604;
wire  [15:0] result3605;
wire  [15:0] result3606;
wire  [15:0] result3607;
wire  [15:0] result3608;
wire  [15:0] result3609;
wire  [15:0] result3610;
wire  [15:0] result3611;
wire  [15:0] result3612;
wire  [15:0] result3613;
wire  [15:0] result3614;
wire  [15:0] result3615;
wire  [15:0] result3616;
wire  [15:0] result3617;
wire  [15:0] result3618;
wire  [15:0] result3619;
wire  [15:0] result3620;
wire  [15:0] result3621;
wire  [15:0] result3622;
wire  [15:0] result3623;
wire  [15:0] result3624;
wire  [15:0] result3625;
wire  [15:0] result3626;
wire  [15:0] result3627;
wire  [15:0] result3628;
wire  [15:0] result3629;
wire  [15:0] result3630;
wire  [15:0] result3631;
wire  [15:0] result3632;
wire  [15:0] result3633;
wire  [15:0] result3634;
wire  [15:0] result3635;
wire  [15:0] result3636;
wire  [15:0] result3637;
wire  [15:0] result3638;
wire  [15:0] result3639;
wire  [15:0] result3640;
wire  [15:0] result3641;
wire  [15:0] result3642;
wire  [15:0] result3643;
wire  [15:0] result3644;
wire  [15:0] result3645;
wire  [15:0] result3646;
wire  [15:0] result3647;
wire  [15:0] result3648;
wire  [15:0] result3649;
wire  [15:0] result3650;
wire  [15:0] result3651;
wire  [15:0] result3652;
wire  [15:0] result3653;
wire  [15:0] result3654;
wire  [15:0] result3655;
wire  [15:0] result3656;
wire  [15:0] result3657;
wire  [15:0] result3658;
wire  [15:0] result3659;
wire  [15:0] result3660;
wire  [15:0] result3661;
wire  [15:0] result3662;
wire  [15:0] result3663;
wire  [15:0] result3664;
wire  [15:0] result3665;
wire  [15:0] result3666;
wire  [15:0] result3667;
wire  [15:0] result3668;
wire  [15:0] result3669;
wire  [15:0] result3670;
wire  [15:0] result3671;
wire  [15:0] result3672;
wire  [15:0] result3673;
wire  [15:0] result3674;
wire  [15:0] result3675;
wire  [15:0] result3676;
wire  [15:0] result3677;
wire  [15:0] result3678;
wire  [15:0] result3679;
wire  [15:0] result3680;
wire  [15:0] result3681;
wire  [15:0] result3682;
wire  [15:0] result3683;
wire  [15:0] result3684;
wire  [15:0] result3685;
wire  [15:0] result3686;
wire  [15:0] result3687;
wire  [15:0] result3688;
wire  [15:0] result3689;
wire  [15:0] result3690;
wire  [15:0] result3691;
wire  [15:0] result3692;
wire  [15:0] result3693;
wire  [15:0] result3694;
wire  [15:0] result3695;
wire  [15:0] result3696;
wire  [15:0] result3697;
wire  [15:0] result3698;
wire  [15:0] result3699;
wire  [15:0] result3700;
wire  [15:0] result3701;
wire  [15:0] result3702;
wire  [15:0] result3703;
wire  [15:0] result3704;
wire  [15:0] result3705;
wire  [15:0] result3706;
wire  [15:0] result3707;
wire  [15:0] result3708;
wire  [15:0] result3709;
wire  [15:0] result3710;
wire  [15:0] result3711;
wire  [15:0] result3712;
wire  [15:0] result3713;
wire  [15:0] result3714;
wire  [15:0] result3715;
wire  [15:0] result3716;
wire  [15:0] result3717;
wire  [15:0] result3718;
wire  [15:0] result3719;
wire  [15:0] result3720;
wire  [15:0] result3721;
wire  [15:0] result3722;
wire  [15:0] result3723;
wire  [15:0] result3724;
wire  [15:0] result3725;
wire  [15:0] result3726;
wire  [15:0] result3727;
wire  [15:0] result3728;
wire  [15:0] result3729;
wire  [15:0] result3730;
wire  [15:0] result3731;
wire  [15:0] result3732;
wire  [15:0] result3733;
wire  [15:0] result3734;
wire  [15:0] result3735;
wire  [15:0] result3736;
wire  [15:0] result3737;
wire  [15:0] result3738;
wire  [15:0] result3739;
wire  [15:0] result3740;
wire  [15:0] result3741;
wire  [15:0] result3742;
wire  [15:0] result3743;
wire  [15:0] result3744;
wire  [15:0] result3745;
wire  [15:0] result3746;
wire  [15:0] result3747;
wire  [15:0] result3748;
wire  [15:0] result3749;
wire  [15:0] result3750;
wire  [15:0] result3751;
wire  [15:0] result3752;
wire  [15:0] result3753;
wire  [15:0] result3754;
wire  [15:0] result3755;
wire  [15:0] result3756;
wire  [15:0] result3757;
wire  [15:0] result3758;
wire  [15:0] result3759;
wire  [15:0] result3760;
wire  [15:0] result3761;
wire  [15:0] result3762;
wire  [15:0] result3763;
wire  [15:0] result3764;
wire  [15:0] result3765;
wire  [15:0] result3766;
wire  [15:0] result3767;
wire  [15:0] result3768;
wire  [15:0] result3769;
wire  [15:0] result3770;
wire  [15:0] result3771;
wire  [15:0] result3772;
wire  [15:0] result3773;
wire  [15:0] result3774;
wire  [15:0] result3775;
wire  [15:0] result3776;
wire  [15:0] result3777;
wire  [15:0] result3778;
wire  [15:0] result3779;
wire  [15:0] result3780;
wire  [15:0] result3781;
wire  [15:0] result3782;
wire  [15:0] result3783;
wire  [15:0] result3784;
wire  [15:0] result3785;
wire  [15:0] result3786;
wire  [15:0] result3787;
wire  [15:0] result3788;
wire  [15:0] result3789;
wire  [15:0] result3790;
wire  [15:0] result3791;
wire  [15:0] result3792;
wire  [15:0] result3793;
wire  [15:0] result3794;
wire  [15:0] result3795;
wire  [15:0] result3796;
wire  [15:0] result3797;
wire  [15:0] result3798;
wire  [15:0] result3799;
wire  [15:0] result3800;
wire  [15:0] result3801;
wire  [15:0] result3802;
wire  [15:0] result3803;
wire  [15:0] result3804;
wire  [15:0] result3805;
wire  [15:0] result3806;
wire  [15:0] result3807;
wire  [15:0] result3808;
wire  [15:0] result3809;
wire  [15:0] result3810;
wire  [15:0] result3811;
wire  [15:0] result3812;
wire  [15:0] result3813;
wire  [15:0] result3814;
wire  [15:0] result3815;
wire  [15:0] result3816;
wire  [15:0] result3817;
wire  [15:0] result3818;
wire  [15:0] result3819;
wire  [15:0] result3820;
wire  [15:0] result3821;
wire  [15:0] result3822;
wire  [15:0] result3823;
wire  [15:0] result3824;
wire  [15:0] result3825;
wire  [15:0] result3826;
wire  [15:0] result3827;
wire  [15:0] result3828;
wire  [15:0] result3829;
wire  [15:0] result3830;
wire  [15:0] result3831;
wire  [15:0] result3832;
wire  [15:0] result3833;
wire  [15:0] result3834;
wire  [15:0] result3835;
wire  [15:0] result3836;
wire  [15:0] result3837;
wire  [15:0] result3838;
wire  [15:0] result3839;
wire  [15:0] result3840;
wire  [15:0] result3841;
wire  [15:0] result3842;
wire  [15:0] result3843;
wire  [15:0] result3844;
wire  [15:0] result3845;
wire  [15:0] result3846;
wire  [15:0] result3847;
wire  [15:0] result3848;
wire  [15:0] result3849;
wire  [15:0] result3850;
wire  [15:0] result3851;
wire  [15:0] result3852;
wire  [15:0] result3853;
wire  [15:0] result3854;
wire  [15:0] result3855;
wire  [15:0] result3856;
wire  [15:0] result3857;
wire  [15:0] result3858;
wire  [15:0] result3859;
wire  [15:0] result3860;
wire  [15:0] result3861;
wire  [15:0] result3862;
wire  [15:0] result3863;
wire  [15:0] result3864;
wire  [15:0] result3865;
wire  [15:0] result3866;
wire  [15:0] result3867;
wire  [15:0] result3868;
wire  [15:0] result3869;
wire  [15:0] result3870;
wire  [15:0] result3871;
wire  [15:0] result3872;
wire  [15:0] result3873;
wire  [15:0] result3874;
wire  [15:0] result3875;
wire  [15:0] result3876;
wire  [15:0] result3877;
wire  [15:0] result3878;
wire  [15:0] result3879;
wire  [15:0] result3880;
wire  [15:0] result3881;
wire  [15:0] result3882;
wire  [15:0] result3883;
wire  [15:0] result3884;
wire  [15:0] result3885;
wire  [15:0] result3886;
wire  [15:0] result3887;
wire  [15:0] result3888;
wire  [15:0] result3889;
wire  [15:0] result3890;
wire  [15:0] result3891;
wire  [15:0] result3892;
wire  [15:0] result3893;
wire  [15:0] result3894;
wire  [15:0] result3895;
wire  [15:0] result3896;
wire  [15:0] result3897;
wire  [15:0] result3898;
wire  [15:0] result3899;
wire  [15:0] result3900;
wire  [15:0] result3901;
wire  [15:0] result3902;
wire  [15:0] result3903;
wire  [15:0] result3904;
wire  [15:0] result3905;
wire  [15:0] result3906;
wire  [15:0] result3907;
wire  [15:0] result3908;
wire  [15:0] result3909;
wire  [15:0] result3910;
wire  [15:0] result3911;
wire  [15:0] result3912;
wire  [15:0] result3913;
wire  [15:0] result3914;
wire  [15:0] result3915;
wire  [15:0] result3916;
wire  [15:0] result3917;
wire  [15:0] result3918;
wire  [15:0] result3919;
wire  [15:0] result3920;
wire  [15:0] result3921;
wire  [15:0] result3922;
wire  [15:0] result3923;
wire  [15:0] result3924;
wire  [15:0] result3925;
wire  [15:0] result3926;
wire  [15:0] result3927;
wire  [15:0] result3928;
wire  [15:0] result3929;
wire  [15:0] result3930;
wire  [15:0] result3931;
wire  [15:0] result3932;
wire  [15:0] result3933;
wire  [15:0] result3934;
wire  [15:0] result3935;
wire  [15:0] result3936;
wire  [15:0] result3937;
wire  [15:0] result3938;
wire  [15:0] result3939;
wire  [15:0] result3940;
wire  [15:0] result3941;
wire  [15:0] result3942;
wire  [15:0] result3943;
wire  [15:0] result3944;
wire  [15:0] result3945;
wire  [15:0] result3946;
wire  [15:0] result3947;
wire  [15:0] result3948;
wire  [15:0] result3949;
wire  [15:0] result3950;
wire  [15:0] result3951;
wire  [15:0] result3952;
wire  [15:0] result3953;
wire  [15:0] result3954;
wire  [15:0] result3955;
wire  [15:0] result3956;
wire  [15:0] result3957;
wire  [15:0] result3958;
wire  [15:0] result3959;
wire  [15:0] result3960;
wire  [15:0] result3961;
wire  [15:0] result3962;
wire  [15:0] result3963;
wire  [15:0] result3964;
wire  [15:0] result3965;
wire  [15:0] result3966;
wire  [15:0] result3967;
wire  [15:0] result3968;
wire  [15:0] result3969;
wire  [15:0] result3970;
wire  [15:0] result3971;
wire  [15:0] result3972;
wire  [15:0] result3973;
wire  [15:0] result3974;
wire  [15:0] result3975;
wire  [15:0] result3976;
wire  [15:0] result3977;
wire  [15:0] result3978;
wire  [15:0] result3979;
wire  [15:0] result3980;
wire  [15:0] result3981;
wire  [15:0] result3982;
wire  [15:0] result3983;
wire  [15:0] result3984;
wire  [15:0] result3985;
wire  [15:0] result3986;
wire  [15:0] result3987;
wire  [15:0] result3988;
wire  [15:0] result3989;
wire  [15:0] result3990;
wire  [15:0] result3991;
wire  [15:0] result3992;
wire  [15:0] result3993;
wire  [15:0] result3994;
wire  [15:0] result3995;
wire  [15:0] result3996;
wire  [15:0] result3997;
wire  [15:0] result3998;
wire  [15:0] result3999;
wire  [15:0] result4000;
wire  [15:0] result4001;
wire  [15:0] result4002;
wire  [15:0] result4003;
wire  [15:0] result4004;
wire  [15:0] result4005;
wire  [15:0] result4006;
wire  [15:0] result4007;
wire  [15:0] result4008;
wire  [15:0] result4009;
wire  [15:0] result4010;
wire  [15:0] result4011;
wire  [15:0] result4012;
wire  [15:0] result4013;
wire  [15:0] result4014;
wire  [15:0] result4015;
wire  [15:0] result4016;
wire  [15:0] result4017;
wire  [15:0] result4018;
wire  [15:0] result4019;
wire  [15:0] result4020;
wire  [15:0] result4021;
wire  [15:0] result4022;
wire  [15:0] result4023;
wire  [15:0] result4024;
wire  [15:0] result4025;
wire  [15:0] result4026;
wire  [15:0] result4027;
wire  [15:0] result4028;
wire  [15:0] result4029;
wire  [15:0] result4030;
wire  [15:0] result4031;
wire  [15:0] result4032;
wire  [15:0] result4033;
wire  [15:0] result4034;
wire  [15:0] result4035;
wire  [15:0] result4036;
wire  [15:0] result4037;
wire  [15:0] result4038;
wire  [15:0] result4039;
wire  [15:0] result4040;
wire  [15:0] result4041;
wire  [15:0] result4042;
wire  [15:0] result4043;
wire  [15:0] result4044;
wire  [15:0] result4045;
wire  [15:0] result4046;
wire  [15:0] result4047;
wire  [15:0] result4048;
wire  [15:0] result4049;
wire  [15:0] result4050;
wire  [15:0] result4051;
wire  [15:0] result4052;
wire  [15:0] result4053;
wire  [15:0] result4054;
wire  [15:0] result4055;
wire  [15:0] result4056;
wire  [15:0] result4057;
wire  [15:0] result4058;
wire  [15:0] result4059;
wire  [15:0] result4060;
wire  [15:0] result4061;
wire  [15:0] result4062;
wire  [15:0] result4063;
wire  [15:0] result4064;
wire  [15:0] result4065;
wire  [15:0] result4066;
wire  [15:0] result4067;
wire  [15:0] result4068;
wire  [15:0] result4069;
wire  [15:0] result4070;
wire  [15:0] result4071;
wire  [15:0] result4072;
wire  [15:0] result4073;
wire  [15:0] result4074;
wire  [15:0] result4075;
wire  [15:0] result4076;
wire  [15:0] result4077;
wire  [15:0] result4078;
wire  [15:0] result4079;
wire  [15:0] result4080;
wire  [15:0] result4081;
wire  [15:0] result4082;
wire  [15:0] result4083;
wire  [15:0] result4084;
wire  [15:0] result4085;
wire  [15:0] result4086;
wire  [15:0] result4087;
wire  [15:0] result4088;
wire  [15:0] result4089;
wire  [15:0] result4090;
wire  [15:0] result4091;
wire  [15:0] result4092;
wire  [15:0] result4093;
wire  [15:0] result4094;
wire  [15:0] result4095;

PE P0 (inp_n0, inp_w0, clk, rst, out_s0, out_e0, result0);

PE P1(inp_n1, out_e1, clk, rst, out_s1, out_e1, result1);
PE P2(inp_n2, out_e2, clk, rst, out_s2, out_e2, result2);
PE P3(inp_n3, out_e3, clk, rst, out_s3, out_e3, result3);
PE P4(inp_n4, out_e4, clk, rst, out_s4, out_e4, result4);
PE P5(inp_n5, out_e5, clk, rst, out_s5, out_e5, result5);
PE P6(inp_n6, out_e6, clk, rst, out_s6, out_e6, result6);
PE P7(inp_n7, out_e7, clk, rst, out_s7, out_e7, result7);
PE P8(inp_n8, out_e8, clk, rst, out_s8, out_e8, result8);
PE P9(inp_n9, out_e9, clk, rst, out_s9, out_e9, result9);
PE P10(inp_n10, out_e10, clk, rst, out_s10, out_e10, result10);
PE P11(inp_n11, out_e11, clk, rst, out_s11, out_e11, result11);
PE P12(inp_n12, out_e12, clk, rst, out_s12, out_e12, result12);
PE P13(inp_n13, out_e13, clk, rst, out_s13, out_e13, result13);
PE P14(inp_n14, out_e14, clk, rst, out_s14, out_e14, result14);
PE P15(inp_n15, out_e15, clk, rst, out_s15, out_e15, result15);
PE P16(inp_n16, out_e16, clk, rst, out_s16, out_e16, result16);
PE P17(inp_n17, out_e17, clk, rst, out_s17, out_e17, result17);
PE P18(inp_n18, out_e18, clk, rst, out_s18, out_e18, result18);
PE P19(inp_n19, out_e19, clk, rst, out_s19, out_e19, result19);
PE P20(inp_n20, out_e20, clk, rst, out_s20, out_e20, result20);
PE P21(inp_n21, out_e21, clk, rst, out_s21, out_e21, result21);
PE P22(inp_n22, out_e22, clk, rst, out_s22, out_e22, result22);
PE P23(inp_n23, out_e23, clk, rst, out_s23, out_e23, result23);
PE P24(inp_n24, out_e24, clk, rst, out_s24, out_e24, result24);
PE P25(inp_n25, out_e25, clk, rst, out_s25, out_e25, result25);
PE P26(inp_n26, out_e26, clk, rst, out_s26, out_e26, result26);
PE P27(inp_n27, out_e27, clk, rst, out_s27, out_e27, result27);
PE P28(inp_n28, out_e28, clk, rst, out_s28, out_e28, result28);
PE P29(inp_n29, out_e29, clk, rst, out_s29, out_e29, result29);
PE P30(inp_n30, out_e30, clk, rst, out_s30, out_e30, result30);
PE P31(inp_n31, out_e31, clk, rst, out_s31, out_e31, result31);
PE P32(inp_n32, out_e32, clk, rst, out_s32, out_e32, result32);
PE P33(inp_n33, out_e33, clk, rst, out_s33, out_e33, result33);
PE P34(inp_n34, out_e34, clk, rst, out_s34, out_e34, result34);
PE P35(inp_n35, out_e35, clk, rst, out_s35, out_e35, result35);
PE P36(inp_n36, out_e36, clk, rst, out_s36, out_e36, result36);
PE P37(inp_n37, out_e37, clk, rst, out_s37, out_e37, result37);
PE P38(inp_n38, out_e38, clk, rst, out_s38, out_e38, result38);
PE P39(inp_n39, out_e39, clk, rst, out_s39, out_e39, result39);
PE P40(inp_n40, out_e40, clk, rst, out_s40, out_e40, result40);
PE P41(inp_n41, out_e41, clk, rst, out_s41, out_e41, result41);
PE P42(inp_n42, out_e42, clk, rst, out_s42, out_e42, result42);
PE P43(inp_n43, out_e43, clk, rst, out_s43, out_e43, result43);
PE P44(inp_n44, out_e44, clk, rst, out_s44, out_e44, result44);
PE P45(inp_n45, out_e45, clk, rst, out_s45, out_e45, result45);
PE P46(inp_n46, out_e46, clk, rst, out_s46, out_e46, result46);
PE P47(inp_n47, out_e47, clk, rst, out_s47, out_e47, result47);
PE P48(inp_n48, out_e48, clk, rst, out_s48, out_e48, result48);
PE P49(inp_n49, out_e49, clk, rst, out_s49, out_e49, result49);
PE P50(inp_n50, out_e50, clk, rst, out_s50, out_e50, result50);
PE P51(inp_n51, out_e51, clk, rst, out_s51, out_e51, result51);
PE P52(inp_n52, out_e52, clk, rst, out_s52, out_e52, result52);
PE P53(inp_n53, out_e53, clk, rst, out_s53, out_e53, result53);
PE P54(inp_n54, out_e54, clk, rst, out_s54, out_e54, result54);
PE P55(inp_n55, out_e55, clk, rst, out_s55, out_e55, result55);
PE P56(inp_n56, out_e56, clk, rst, out_s56, out_e56, result56);
PE P57(inp_n57, out_e57, clk, rst, out_s57, out_e57, result57);
PE P58(inp_n58, out_e58, clk, rst, out_s58, out_e58, result58);
PE P59(inp_n59, out_e59, clk, rst, out_s59, out_e59, result59);
PE P60(inp_n60, out_e60, clk, rst, out_s60, out_e60, result60);
PE P61(inp_n61, out_e61, clk, rst, out_s61, out_e61, result61);
PE P62(inp_n62, out_e62, clk, rst, out_s62, out_e62, result62);
PE P63(inp_n63, out_e63, clk, rst, out_s63, out_e63, result63);

PE P64(out_s0, inp_w64, clk, rst, out_s64, out_e64, result64);
PE P128(out_s64, inp_w128, clk, rst, out_s128, out_e128, result128);
PE P192(out_s128, inp_w192, clk, rst, out_s192, out_e192, result192);
PE P256(out_s192, inp_w256, clk, rst, out_s256, out_e256, result256);
PE P320(out_s256, inp_w320, clk, rst, out_s320, out_e320, result320);
PE P384(out_s320, inp_w384, clk, rst, out_s384, out_e384, result384);
PE P448(out_s384, inp_w448, clk, rst, out_s448, out_e448, result448);
PE P512(out_s448, inp_w512, clk, rst, out_s512, out_e512, result512);
PE P576(out_s512, inp_w576, clk, rst, out_s576, out_e576, result576);
PE P640(out_s576, inp_w640, clk, rst, out_s640, out_e640, result640);
PE P704(out_s640, inp_w704, clk, rst, out_s704, out_e704, result704);
PE P768(out_s704, inp_w768, clk, rst, out_s768, out_e768, result768);
PE P832(out_s768, inp_w832, clk, rst, out_s832, out_e832, result832);
PE P896(out_s832, inp_w896, clk, rst, out_s896, out_e896, result896);
PE P960(out_s896, inp_w960, clk, rst, out_s960, out_e960, result960);
PE P1024(out_s960, inp_w1024, clk, rst, out_s1024, out_e1024, result1024);
PE P1088(out_s1024, inp_w1088, clk, rst, out_s1088, out_e1088, result1088);
PE P1152(out_s1088, inp_w1152, clk, rst, out_s1152, out_e1152, result1152);
PE P1216(out_s1152, inp_w1216, clk, rst, out_s1216, out_e1216, result1216);
PE P1280(out_s1216, inp_w1280, clk, rst, out_s1280, out_e1280, result1280);
PE P1344(out_s1280, inp_w1344, clk, rst, out_s1344, out_e1344, result1344);
PE P1408(out_s1344, inp_w1408, clk, rst, out_s1408, out_e1408, result1408);
PE P1472(out_s1408, inp_w1472, clk, rst, out_s1472, out_e1472, result1472);
PE P1536(out_s1472, inp_w1536, clk, rst, out_s1536, out_e1536, result1536);
PE P1600(out_s1536, inp_w1600, clk, rst, out_s1600, out_e1600, result1600);
PE P1664(out_s1600, inp_w1664, clk, rst, out_s1664, out_e1664, result1664);
PE P1728(out_s1664, inp_w1728, clk, rst, out_s1728, out_e1728, result1728);
PE P1792(out_s1728, inp_w1792, clk, rst, out_s1792, out_e1792, result1792);
PE P1856(out_s1792, inp_w1856, clk, rst, out_s1856, out_e1856, result1856);
PE P1920(out_s1856, inp_w1920, clk, rst, out_s1920, out_e1920, result1920);
PE P1984(out_s1920, inp_w1984, clk, rst, out_s1984, out_e1984, result1984);
PE P2048(out_s1984, inp_w2048, clk, rst, out_s2048, out_e2048, result2048);
PE P2112(out_s2048, inp_w2112, clk, rst, out_s2112, out_e2112, result2112);
PE P2176(out_s2112, inp_w2176, clk, rst, out_s2176, out_e2176, result2176);
PE P2240(out_s2176, inp_w2240, clk, rst, out_s2240, out_e2240, result2240);
PE P2304(out_s2240, inp_w2304, clk, rst, out_s2304, out_e2304, result2304);
PE P2368(out_s2304, inp_w2368, clk, rst, out_s2368, out_e2368, result2368);
PE P2432(out_s2368, inp_w2432, clk, rst, out_s2432, out_e2432, result2432);
PE P2496(out_s2432, inp_w2496, clk, rst, out_s2496, out_e2496, result2496);
PE P2560(out_s2496, inp_w2560, clk, rst, out_s2560, out_e2560, result2560);
PE P2624(out_s2560, inp_w2624, clk, rst, out_s2624, out_e2624, result2624);
PE P2688(out_s2624, inp_w2688, clk, rst, out_s2688, out_e2688, result2688);
PE P2752(out_s2688, inp_w2752, clk, rst, out_s2752, out_e2752, result2752);
PE P2816(out_s2752, inp_w2816, clk, rst, out_s2816, out_e2816, result2816);
PE P2880(out_s2816, inp_w2880, clk, rst, out_s2880, out_e2880, result2880);
PE P2944(out_s2880, inp_w2944, clk, rst, out_s2944, out_e2944, result2944);
PE P3008(out_s2944, inp_w3008, clk, rst, out_s3008, out_e3008, result3008);
PE P3072(out_s3008, inp_w3072, clk, rst, out_s3072, out_e3072, result3072);
PE P3136(out_s3072, inp_w3136, clk, rst, out_s3136, out_e3136, result3136);
PE P3200(out_s3136, inp_w3200, clk, rst, out_s3200, out_e3200, result3200);
PE P3264(out_s3200, inp_w3264, clk, rst, out_s3264, out_e3264, result3264);
PE P3328(out_s3264, inp_w3328, clk, rst, out_s3328, out_e3328, result3328);
PE P3392(out_s3328, inp_w3392, clk, rst, out_s3392, out_e3392, result3392);
PE P3456(out_s3392, inp_w3456, clk, rst, out_s3456, out_e3456, result3456);
PE P3520(out_s3456, inp_w3520, clk, rst, out_s3520, out_e3520, result3520);
PE P3584(out_s3520, inp_w3584, clk, rst, out_s3584, out_e3584, result3584);
PE P3648(out_s3584, inp_w3648, clk, rst, out_s3648, out_e3648, result3648);
PE P3712(out_s3648, inp_w3712, clk, rst, out_s3712, out_e3712, result3712);
PE P3776(out_s3712, inp_w3776, clk, rst, out_s3776, out_e3776, result3776);
PE P3840(out_s3776, inp_w3840, clk, rst, out_s3840, out_e3840, result3840);
PE P3904(out_s3840, inp_w3904, clk, rst, out_s3904, out_e3904, result3904);
PE P3968(out_s3904, inp_w3968, clk, rst, out_s3968, out_e3968, result3968);
PE P4032(out_s3968, inp_w4032, clk, rst, out_s4032, out_e4032, result4032);

PE P65(out_s1, out_e64, clk, rst, out_s65, out_e65, result65);
PE P66(out_s2, out_e65, clk, rst, out_s66, out_e66, result66);
PE P67(out_s3, out_e66, clk, rst, out_s67, out_e67, result67);
PE P68(out_s4, out_e67, clk, rst, out_s68, out_e68, result68);
PE P69(out_s5, out_e68, clk, rst, out_s69, out_e69, result69);
PE P70(out_s6, out_e69, clk, rst, out_s70, out_e70, result70);
PE P71(out_s7, out_e70, clk, rst, out_s71, out_e71, result71);
PE P72(out_s8, out_e71, clk, rst, out_s72, out_e72, result72);
PE P73(out_s9, out_e72, clk, rst, out_s73, out_e73, result73);
PE P74(out_s10, out_e73, clk, rst, out_s74, out_e74, result74);
PE P75(out_s11, out_e74, clk, rst, out_s75, out_e75, result75);
PE P76(out_s12, out_e75, clk, rst, out_s76, out_e76, result76);
PE P77(out_s13, out_e76, clk, rst, out_s77, out_e77, result77);
PE P78(out_s14, out_e77, clk, rst, out_s78, out_e78, result78);
PE P79(out_s15, out_e78, clk, rst, out_s79, out_e79, result79);
PE P80(out_s16, out_e79, clk, rst, out_s80, out_e80, result80);
PE P81(out_s17, out_e80, clk, rst, out_s81, out_e81, result81);
PE P82(out_s18, out_e81, clk, rst, out_s82, out_e82, result82);
PE P83(out_s19, out_e82, clk, rst, out_s83, out_e83, result83);
PE P84(out_s20, out_e83, clk, rst, out_s84, out_e84, result84);
PE P85(out_s21, out_e84, clk, rst, out_s85, out_e85, result85);
PE P86(out_s22, out_e85, clk, rst, out_s86, out_e86, result86);
PE P87(out_s23, out_e86, clk, rst, out_s87, out_e87, result87);
PE P88(out_s24, out_e87, clk, rst, out_s88, out_e88, result88);
PE P89(out_s25, out_e88, clk, rst, out_s89, out_e89, result89);
PE P90(out_s26, out_e89, clk, rst, out_s90, out_e90, result90);
PE P91(out_s27, out_e90, clk, rst, out_s91, out_e91, result91);
PE P92(out_s28, out_e91, clk, rst, out_s92, out_e92, result92);
PE P93(out_s29, out_e92, clk, rst, out_s93, out_e93, result93);
PE P94(out_s30, out_e93, clk, rst, out_s94, out_e94, result94);
PE P95(out_s31, out_e94, clk, rst, out_s95, out_e95, result95);
PE P96(out_s32, out_e95, clk, rst, out_s96, out_e96, result96);
PE P97(out_s33, out_e96, clk, rst, out_s97, out_e97, result97);
PE P98(out_s34, out_e97, clk, rst, out_s98, out_e98, result98);
PE P99(out_s35, out_e98, clk, rst, out_s99, out_e99, result99);
PE P100(out_s36, out_e99, clk, rst, out_s100, out_e100, result100);
PE P101(out_s37, out_e100, clk, rst, out_s101, out_e101, result101);
PE P102(out_s38, out_e101, clk, rst, out_s102, out_e102, result102);
PE P103(out_s39, out_e102, clk, rst, out_s103, out_e103, result103);
PE P104(out_s40, out_e103, clk, rst, out_s104, out_e104, result104);
PE P105(out_s41, out_e104, clk, rst, out_s105, out_e105, result105);
PE P106(out_s42, out_e105, clk, rst, out_s106, out_e106, result106);
PE P107(out_s43, out_e106, clk, rst, out_s107, out_e107, result107);
PE P108(out_s44, out_e107, clk, rst, out_s108, out_e108, result108);
PE P109(out_s45, out_e108, clk, rst, out_s109, out_e109, result109);
PE P110(out_s46, out_e109, clk, rst, out_s110, out_e110, result110);
PE P111(out_s47, out_e110, clk, rst, out_s111, out_e111, result111);
PE P112(out_s48, out_e111, clk, rst, out_s112, out_e112, result112);
PE P113(out_s49, out_e112, clk, rst, out_s113, out_e113, result113);
PE P114(out_s50, out_e113, clk, rst, out_s114, out_e114, result114);
PE P115(out_s51, out_e114, clk, rst, out_s115, out_e115, result115);
PE P116(out_s52, out_e115, clk, rst, out_s116, out_e116, result116);
PE P117(out_s53, out_e116, clk, rst, out_s117, out_e117, result117);
PE P118(out_s54, out_e117, clk, rst, out_s118, out_e118, result118);
PE P119(out_s55, out_e118, clk, rst, out_s119, out_e119, result119);
PE P120(out_s56, out_e119, clk, rst, out_s120, out_e120, result120);
PE P121(out_s57, out_e120, clk, rst, out_s121, out_e121, result121);
PE P122(out_s58, out_e121, clk, rst, out_s122, out_e122, result122);
PE P123(out_s59, out_e122, clk, rst, out_s123, out_e123, result123);
PE P124(out_s60, out_e123, clk, rst, out_s124, out_e124, result124);
PE P125(out_s61, out_e124, clk, rst, out_s125, out_e125, result125);
PE P126(out_s62, out_e125, clk, rst, out_s126, out_e126, result126);
PE P127(out_s63, out_e126, clk, rst, out_s127, out_e127, result127);

PE P129(out_s65, out_e128, clk, rst, out_s129, out_e129, result129);
PE P130(out_s66, out_e129, clk, rst, out_s130, out_e130, result130);
PE P131(out_s67, out_e130, clk, rst, out_s131, out_e131, result131);
PE P132(out_s68, out_e131, clk, rst, out_s132, out_e132, result132);
PE P133(out_s69, out_e132, clk, rst, out_s133, out_e133, result133);
PE P134(out_s70, out_e133, clk, rst, out_s134, out_e134, result134);
PE P135(out_s71, out_e134, clk, rst, out_s135, out_e135, result135);
PE P136(out_s72, out_e135, clk, rst, out_s136, out_e136, result136);
PE P137(out_s73, out_e136, clk, rst, out_s137, out_e137, result137);
PE P138(out_s74, out_e137, clk, rst, out_s138, out_e138, result138);
PE P139(out_s75, out_e138, clk, rst, out_s139, out_e139, result139);
PE P140(out_s76, out_e139, clk, rst, out_s140, out_e140, result140);
PE P141(out_s77, out_e140, clk, rst, out_s141, out_e141, result141);
PE P142(out_s78, out_e141, clk, rst, out_s142, out_e142, result142);
PE P143(out_s79, out_e142, clk, rst, out_s143, out_e143, result143);
PE P144(out_s80, out_e143, clk, rst, out_s144, out_e144, result144);
PE P145(out_s81, out_e144, clk, rst, out_s145, out_e145, result145);
PE P146(out_s82, out_e145, clk, rst, out_s146, out_e146, result146);
PE P147(out_s83, out_e146, clk, rst, out_s147, out_e147, result147);
PE P148(out_s84, out_e147, clk, rst, out_s148, out_e148, result148);
PE P149(out_s85, out_e148, clk, rst, out_s149, out_e149, result149);
PE P150(out_s86, out_e149, clk, rst, out_s150, out_e150, result150);
PE P151(out_s87, out_e150, clk, rst, out_s151, out_e151, result151);
PE P152(out_s88, out_e151, clk, rst, out_s152, out_e152, result152);
PE P153(out_s89, out_e152, clk, rst, out_s153, out_e153, result153);
PE P154(out_s90, out_e153, clk, rst, out_s154, out_e154, result154);
PE P155(out_s91, out_e154, clk, rst, out_s155, out_e155, result155);
PE P156(out_s92, out_e155, clk, rst, out_s156, out_e156, result156);
PE P157(out_s93, out_e156, clk, rst, out_s157, out_e157, result157);
PE P158(out_s94, out_e157, clk, rst, out_s158, out_e158, result158);
PE P159(out_s95, out_e158, clk, rst, out_s159, out_e159, result159);
PE P160(out_s96, out_e159, clk, rst, out_s160, out_e160, result160);
PE P161(out_s97, out_e160, clk, rst, out_s161, out_e161, result161);
PE P162(out_s98, out_e161, clk, rst, out_s162, out_e162, result162);
PE P163(out_s99, out_e162, clk, rst, out_s163, out_e163, result163);
PE P164(out_s100, out_e163, clk, rst, out_s164, out_e164, result164);
PE P165(out_s101, out_e164, clk, rst, out_s165, out_e165, result165);
PE P166(out_s102, out_e165, clk, rst, out_s166, out_e166, result166);
PE P167(out_s103, out_e166, clk, rst, out_s167, out_e167, result167);
PE P168(out_s104, out_e167, clk, rst, out_s168, out_e168, result168);
PE P169(out_s105, out_e168, clk, rst, out_s169, out_e169, result169);
PE P170(out_s106, out_e169, clk, rst, out_s170, out_e170, result170);
PE P171(out_s107, out_e170, clk, rst, out_s171, out_e171, result171);
PE P172(out_s108, out_e171, clk, rst, out_s172, out_e172, result172);
PE P173(out_s109, out_e172, clk, rst, out_s173, out_e173, result173);
PE P174(out_s110, out_e173, clk, rst, out_s174, out_e174, result174);
PE P175(out_s111, out_e174, clk, rst, out_s175, out_e175, result175);
PE P176(out_s112, out_e175, clk, rst, out_s176, out_e176, result176);
PE P177(out_s113, out_e176, clk, rst, out_s177, out_e177, result177);
PE P178(out_s114, out_e177, clk, rst, out_s178, out_e178, result178);
PE P179(out_s115, out_e178, clk, rst, out_s179, out_e179, result179);
PE P180(out_s116, out_e179, clk, rst, out_s180, out_e180, result180);
PE P181(out_s117, out_e180, clk, rst, out_s181, out_e181, result181);
PE P182(out_s118, out_e181, clk, rst, out_s182, out_e182, result182);
PE P183(out_s119, out_e182, clk, rst, out_s183, out_e183, result183);
PE P184(out_s120, out_e183, clk, rst, out_s184, out_e184, result184);
PE P185(out_s121, out_e184, clk, rst, out_s185, out_e185, result185);
PE P186(out_s122, out_e185, clk, rst, out_s186, out_e186, result186);
PE P187(out_s123, out_e186, clk, rst, out_s187, out_e187, result187);
PE P188(out_s124, out_e187, clk, rst, out_s188, out_e188, result188);
PE P189(out_s125, out_e188, clk, rst, out_s189, out_e189, result189);
PE P190(out_s126, out_e189, clk, rst, out_s190, out_e190, result190);
PE P191(out_s127, out_e190, clk, rst, out_s191, out_e191, result191);

PE P193(out_s129, out_e192, clk, rst, out_s193, out_e193, result193);
PE P194(out_s130, out_e193, clk, rst, out_s194, out_e194, result194);
PE P195(out_s131, out_e194, clk, rst, out_s195, out_e195, result195);
PE P196(out_s132, out_e195, clk, rst, out_s196, out_e196, result196);
PE P197(out_s133, out_e196, clk, rst, out_s197, out_e197, result197);
PE P198(out_s134, out_e197, clk, rst, out_s198, out_e198, result198);
PE P199(out_s135, out_e198, clk, rst, out_s199, out_e199, result199);
PE P200(out_s136, out_e199, clk, rst, out_s200, out_e200, result200);
PE P201(out_s137, out_e200, clk, rst, out_s201, out_e201, result201);
PE P202(out_s138, out_e201, clk, rst, out_s202, out_e202, result202);
PE P203(out_s139, out_e202, clk, rst, out_s203, out_e203, result203);
PE P204(out_s140, out_e203, clk, rst, out_s204, out_e204, result204);
PE P205(out_s141, out_e204, clk, rst, out_s205, out_e205, result205);
PE P206(out_s142, out_e205, clk, rst, out_s206, out_e206, result206);
PE P207(out_s143, out_e206, clk, rst, out_s207, out_e207, result207);
PE P208(out_s144, out_e207, clk, rst, out_s208, out_e208, result208);
PE P209(out_s145, out_e208, clk, rst, out_s209, out_e209, result209);
PE P210(out_s146, out_e209, clk, rst, out_s210, out_e210, result210);
PE P211(out_s147, out_e210, clk, rst, out_s211, out_e211, result211);
PE P212(out_s148, out_e211, clk, rst, out_s212, out_e212, result212);
PE P213(out_s149, out_e212, clk, rst, out_s213, out_e213, result213);
PE P214(out_s150, out_e213, clk, rst, out_s214, out_e214, result214);
PE P215(out_s151, out_e214, clk, rst, out_s215, out_e215, result215);
PE P216(out_s152, out_e215, clk, rst, out_s216, out_e216, result216);
PE P217(out_s153, out_e216, clk, rst, out_s217, out_e217, result217);
PE P218(out_s154, out_e217, clk, rst, out_s218, out_e218, result218);
PE P219(out_s155, out_e218, clk, rst, out_s219, out_e219, result219);
PE P220(out_s156, out_e219, clk, rst, out_s220, out_e220, result220);
PE P221(out_s157, out_e220, clk, rst, out_s221, out_e221, result221);
PE P222(out_s158, out_e221, clk, rst, out_s222, out_e222, result222);
PE P223(out_s159, out_e222, clk, rst, out_s223, out_e223, result223);
PE P224(out_s160, out_e223, clk, rst, out_s224, out_e224, result224);
PE P225(out_s161, out_e224, clk, rst, out_s225, out_e225, result225);
PE P226(out_s162, out_e225, clk, rst, out_s226, out_e226, result226);
PE P227(out_s163, out_e226, clk, rst, out_s227, out_e227, result227);
PE P228(out_s164, out_e227, clk, rst, out_s228, out_e228, result228);
PE P229(out_s165, out_e228, clk, rst, out_s229, out_e229, result229);
PE P230(out_s166, out_e229, clk, rst, out_s230, out_e230, result230);
PE P231(out_s167, out_e230, clk, rst, out_s231, out_e231, result231);
PE P232(out_s168, out_e231, clk, rst, out_s232, out_e232, result232);
PE P233(out_s169, out_e232, clk, rst, out_s233, out_e233, result233);
PE P234(out_s170, out_e233, clk, rst, out_s234, out_e234, result234);
PE P235(out_s171, out_e234, clk, rst, out_s235, out_e235, result235);
PE P236(out_s172, out_e235, clk, rst, out_s236, out_e236, result236);
PE P237(out_s173, out_e236, clk, rst, out_s237, out_e237, result237);
PE P238(out_s174, out_e237, clk, rst, out_s238, out_e238, result238);
PE P239(out_s175, out_e238, clk, rst, out_s239, out_e239, result239);
PE P240(out_s176, out_e239, clk, rst, out_s240, out_e240, result240);
PE P241(out_s177, out_e240, clk, rst, out_s241, out_e241, result241);
PE P242(out_s178, out_e241, clk, rst, out_s242, out_e242, result242);
PE P243(out_s179, out_e242, clk, rst, out_s243, out_e243, result243);
PE P244(out_s180, out_e243, clk, rst, out_s244, out_e244, result244);
PE P245(out_s181, out_e244, clk, rst, out_s245, out_e245, result245);
PE P246(out_s182, out_e245, clk, rst, out_s246, out_e246, result246);
PE P247(out_s183, out_e246, clk, rst, out_s247, out_e247, result247);
PE P248(out_s184, out_e247, clk, rst, out_s248, out_e248, result248);
PE P249(out_s185, out_e248, clk, rst, out_s249, out_e249, result249);
PE P250(out_s186, out_e249, clk, rst, out_s250, out_e250, result250);
PE P251(out_s187, out_e250, clk, rst, out_s251, out_e251, result251);
PE P252(out_s188, out_e251, clk, rst, out_s252, out_e252, result252);
PE P253(out_s189, out_e252, clk, rst, out_s253, out_e253, result253);
PE P254(out_s190, out_e253, clk, rst, out_s254, out_e254, result254);
PE P255(out_s191, out_e254, clk, rst, out_s255, out_e255, result255);

PE P257(out_s193, out_e256, clk, rst, out_s257, out_e257, result257);
PE P258(out_s194, out_e257, clk, rst, out_s258, out_e258, result258);
PE P259(out_s195, out_e258, clk, rst, out_s259, out_e259, result259);
PE P260(out_s196, out_e259, clk, rst, out_s260, out_e260, result260);
PE P261(out_s197, out_e260, clk, rst, out_s261, out_e261, result261);
PE P262(out_s198, out_e261, clk, rst, out_s262, out_e262, result262);
PE P263(out_s199, out_e262, clk, rst, out_s263, out_e263, result263);
PE P264(out_s200, out_e263, clk, rst, out_s264, out_e264, result264);
PE P265(out_s201, out_e264, clk, rst, out_s265, out_e265, result265);
PE P266(out_s202, out_e265, clk, rst, out_s266, out_e266, result266);
PE P267(out_s203, out_e266, clk, rst, out_s267, out_e267, result267);
PE P268(out_s204, out_e267, clk, rst, out_s268, out_e268, result268);
PE P269(out_s205, out_e268, clk, rst, out_s269, out_e269, result269);
PE P270(out_s206, out_e269, clk, rst, out_s270, out_e270, result270);
PE P271(out_s207, out_e270, clk, rst, out_s271, out_e271, result271);
PE P272(out_s208, out_e271, clk, rst, out_s272, out_e272, result272);
PE P273(out_s209, out_e272, clk, rst, out_s273, out_e273, result273);
PE P274(out_s210, out_e273, clk, rst, out_s274, out_e274, result274);
PE P275(out_s211, out_e274, clk, rst, out_s275, out_e275, result275);
PE P276(out_s212, out_e275, clk, rst, out_s276, out_e276, result276);
PE P277(out_s213, out_e276, clk, rst, out_s277, out_e277, result277);
PE P278(out_s214, out_e277, clk, rst, out_s278, out_e278, result278);
PE P279(out_s215, out_e278, clk, rst, out_s279, out_e279, result279);
PE P280(out_s216, out_e279, clk, rst, out_s280, out_e280, result280);
PE P281(out_s217, out_e280, clk, rst, out_s281, out_e281, result281);
PE P282(out_s218, out_e281, clk, rst, out_s282, out_e282, result282);
PE P283(out_s219, out_e282, clk, rst, out_s283, out_e283, result283);
PE P284(out_s220, out_e283, clk, rst, out_s284, out_e284, result284);
PE P285(out_s221, out_e284, clk, rst, out_s285, out_e285, result285);
PE P286(out_s222, out_e285, clk, rst, out_s286, out_e286, result286);
PE P287(out_s223, out_e286, clk, rst, out_s287, out_e287, result287);
PE P288(out_s224, out_e287, clk, rst, out_s288, out_e288, result288);
PE P289(out_s225, out_e288, clk, rst, out_s289, out_e289, result289);
PE P290(out_s226, out_e289, clk, rst, out_s290, out_e290, result290);
PE P291(out_s227, out_e290, clk, rst, out_s291, out_e291, result291);
PE P292(out_s228, out_e291, clk, rst, out_s292, out_e292, result292);
PE P293(out_s229, out_e292, clk, rst, out_s293, out_e293, result293);
PE P294(out_s230, out_e293, clk, rst, out_s294, out_e294, result294);
PE P295(out_s231, out_e294, clk, rst, out_s295, out_e295, result295);
PE P296(out_s232, out_e295, clk, rst, out_s296, out_e296, result296);
PE P297(out_s233, out_e296, clk, rst, out_s297, out_e297, result297);
PE P298(out_s234, out_e297, clk, rst, out_s298, out_e298, result298);
PE P299(out_s235, out_e298, clk, rst, out_s299, out_e299, result299);
PE P300(out_s236, out_e299, clk, rst, out_s300, out_e300, result300);
PE P301(out_s237, out_e300, clk, rst, out_s301, out_e301, result301);
PE P302(out_s238, out_e301, clk, rst, out_s302, out_e302, result302);
PE P303(out_s239, out_e302, clk, rst, out_s303, out_e303, result303);
PE P304(out_s240, out_e303, clk, rst, out_s304, out_e304, result304);
PE P305(out_s241, out_e304, clk, rst, out_s305, out_e305, result305);
PE P306(out_s242, out_e305, clk, rst, out_s306, out_e306, result306);
PE P307(out_s243, out_e306, clk, rst, out_s307, out_e307, result307);
PE P308(out_s244, out_e307, clk, rst, out_s308, out_e308, result308);
PE P309(out_s245, out_e308, clk, rst, out_s309, out_e309, result309);
PE P310(out_s246, out_e309, clk, rst, out_s310, out_e310, result310);
PE P311(out_s247, out_e310, clk, rst, out_s311, out_e311, result311);
PE P312(out_s248, out_e311, clk, rst, out_s312, out_e312, result312);
PE P313(out_s249, out_e312, clk, rst, out_s313, out_e313, result313);
PE P314(out_s250, out_e313, clk, rst, out_s314, out_e314, result314);
PE P315(out_s251, out_e314, clk, rst, out_s315, out_e315, result315);
PE P316(out_s252, out_e315, clk, rst, out_s316, out_e316, result316);
PE P317(out_s253, out_e316, clk, rst, out_s317, out_e317, result317);
PE P318(out_s254, out_e317, clk, rst, out_s318, out_e318, result318);
PE P319(out_s255, out_e318, clk, rst, out_s319, out_e319, result319);

PE P321(out_s257, out_e320, clk, rst, out_s321, out_e321, result321);
PE P322(out_s258, out_e321, clk, rst, out_s322, out_e322, result322);
PE P323(out_s259, out_e322, clk, rst, out_s323, out_e323, result323);
PE P324(out_s260, out_e323, clk, rst, out_s324, out_e324, result324);
PE P325(out_s261, out_e324, clk, rst, out_s325, out_e325, result325);
PE P326(out_s262, out_e325, clk, rst, out_s326, out_e326, result326);
PE P327(out_s263, out_e326, clk, rst, out_s327, out_e327, result327);
PE P328(out_s264, out_e327, clk, rst, out_s328, out_e328, result328);
PE P329(out_s265, out_e328, clk, rst, out_s329, out_e329, result329);
PE P330(out_s266, out_e329, clk, rst, out_s330, out_e330, result330);
PE P331(out_s267, out_e330, clk, rst, out_s331, out_e331, result331);
PE P332(out_s268, out_e331, clk, rst, out_s332, out_e332, result332);
PE P333(out_s269, out_e332, clk, rst, out_s333, out_e333, result333);
PE P334(out_s270, out_e333, clk, rst, out_s334, out_e334, result334);
PE P335(out_s271, out_e334, clk, rst, out_s335, out_e335, result335);
PE P336(out_s272, out_e335, clk, rst, out_s336, out_e336, result336);
PE P337(out_s273, out_e336, clk, rst, out_s337, out_e337, result337);
PE P338(out_s274, out_e337, clk, rst, out_s338, out_e338, result338);
PE P339(out_s275, out_e338, clk, rst, out_s339, out_e339, result339);
PE P340(out_s276, out_e339, clk, rst, out_s340, out_e340, result340);
PE P341(out_s277, out_e340, clk, rst, out_s341, out_e341, result341);
PE P342(out_s278, out_e341, clk, rst, out_s342, out_e342, result342);
PE P343(out_s279, out_e342, clk, rst, out_s343, out_e343, result343);
PE P344(out_s280, out_e343, clk, rst, out_s344, out_e344, result344);
PE P345(out_s281, out_e344, clk, rst, out_s345, out_e345, result345);
PE P346(out_s282, out_e345, clk, rst, out_s346, out_e346, result346);
PE P347(out_s283, out_e346, clk, rst, out_s347, out_e347, result347);
PE P348(out_s284, out_e347, clk, rst, out_s348, out_e348, result348);
PE P349(out_s285, out_e348, clk, rst, out_s349, out_e349, result349);
PE P350(out_s286, out_e349, clk, rst, out_s350, out_e350, result350);
PE P351(out_s287, out_e350, clk, rst, out_s351, out_e351, result351);
PE P352(out_s288, out_e351, clk, rst, out_s352, out_e352, result352);
PE P353(out_s289, out_e352, clk, rst, out_s353, out_e353, result353);
PE P354(out_s290, out_e353, clk, rst, out_s354, out_e354, result354);
PE P355(out_s291, out_e354, clk, rst, out_s355, out_e355, result355);
PE P356(out_s292, out_e355, clk, rst, out_s356, out_e356, result356);
PE P357(out_s293, out_e356, clk, rst, out_s357, out_e357, result357);
PE P358(out_s294, out_e357, clk, rst, out_s358, out_e358, result358);
PE P359(out_s295, out_e358, clk, rst, out_s359, out_e359, result359);
PE P360(out_s296, out_e359, clk, rst, out_s360, out_e360, result360);
PE P361(out_s297, out_e360, clk, rst, out_s361, out_e361, result361);
PE P362(out_s298, out_e361, clk, rst, out_s362, out_e362, result362);
PE P363(out_s299, out_e362, clk, rst, out_s363, out_e363, result363);
PE P364(out_s300, out_e363, clk, rst, out_s364, out_e364, result364);
PE P365(out_s301, out_e364, clk, rst, out_s365, out_e365, result365);
PE P366(out_s302, out_e365, clk, rst, out_s366, out_e366, result366);
PE P367(out_s303, out_e366, clk, rst, out_s367, out_e367, result367);
PE P368(out_s304, out_e367, clk, rst, out_s368, out_e368, result368);
PE P369(out_s305, out_e368, clk, rst, out_s369, out_e369, result369);
PE P370(out_s306, out_e369, clk, rst, out_s370, out_e370, result370);
PE P371(out_s307, out_e370, clk, rst, out_s371, out_e371, result371);
PE P372(out_s308, out_e371, clk, rst, out_s372, out_e372, result372);
PE P373(out_s309, out_e372, clk, rst, out_s373, out_e373, result373);
PE P374(out_s310, out_e373, clk, rst, out_s374, out_e374, result374);
PE P375(out_s311, out_e374, clk, rst, out_s375, out_e375, result375);
PE P376(out_s312, out_e375, clk, rst, out_s376, out_e376, result376);
PE P377(out_s313, out_e376, clk, rst, out_s377, out_e377, result377);
PE P378(out_s314, out_e377, clk, rst, out_s378, out_e378, result378);
PE P379(out_s315, out_e378, clk, rst, out_s379, out_e379, result379);
PE P380(out_s316, out_e379, clk, rst, out_s380, out_e380, result380);
PE P381(out_s317, out_e380, clk, rst, out_s381, out_e381, result381);
PE P382(out_s318, out_e381, clk, rst, out_s382, out_e382, result382);
PE P383(out_s319, out_e382, clk, rst, out_s383, out_e383, result383);

PE P385(out_s321, out_e384, clk, rst, out_s385, out_e385, result385);
PE P386(out_s322, out_e385, clk, rst, out_s386, out_e386, result386);
PE P387(out_s323, out_e386, clk, rst, out_s387, out_e387, result387);
PE P388(out_s324, out_e387, clk, rst, out_s388, out_e388, result388);
PE P389(out_s325, out_e388, clk, rst, out_s389, out_e389, result389);
PE P390(out_s326, out_e389, clk, rst, out_s390, out_e390, result390);
PE P391(out_s327, out_e390, clk, rst, out_s391, out_e391, result391);
PE P392(out_s328, out_e391, clk, rst, out_s392, out_e392, result392);
PE P393(out_s329, out_e392, clk, rst, out_s393, out_e393, result393);
PE P394(out_s330, out_e393, clk, rst, out_s394, out_e394, result394);
PE P395(out_s331, out_e394, clk, rst, out_s395, out_e395, result395);
PE P396(out_s332, out_e395, clk, rst, out_s396, out_e396, result396);
PE P397(out_s333, out_e396, clk, rst, out_s397, out_e397, result397);
PE P398(out_s334, out_e397, clk, rst, out_s398, out_e398, result398);
PE P399(out_s335, out_e398, clk, rst, out_s399, out_e399, result399);
PE P400(out_s336, out_e399, clk, rst, out_s400, out_e400, result400);
PE P401(out_s337, out_e400, clk, rst, out_s401, out_e401, result401);
PE P402(out_s338, out_e401, clk, rst, out_s402, out_e402, result402);
PE P403(out_s339, out_e402, clk, rst, out_s403, out_e403, result403);
PE P404(out_s340, out_e403, clk, rst, out_s404, out_e404, result404);
PE P405(out_s341, out_e404, clk, rst, out_s405, out_e405, result405);
PE P406(out_s342, out_e405, clk, rst, out_s406, out_e406, result406);
PE P407(out_s343, out_e406, clk, rst, out_s407, out_e407, result407);
PE P408(out_s344, out_e407, clk, rst, out_s408, out_e408, result408);
PE P409(out_s345, out_e408, clk, rst, out_s409, out_e409, result409);
PE P410(out_s346, out_e409, clk, rst, out_s410, out_e410, result410);
PE P411(out_s347, out_e410, clk, rst, out_s411, out_e411, result411);
PE P412(out_s348, out_e411, clk, rst, out_s412, out_e412, result412);
PE P413(out_s349, out_e412, clk, rst, out_s413, out_e413, result413);
PE P414(out_s350, out_e413, clk, rst, out_s414, out_e414, result414);
PE P415(out_s351, out_e414, clk, rst, out_s415, out_e415, result415);
PE P416(out_s352, out_e415, clk, rst, out_s416, out_e416, result416);
PE P417(out_s353, out_e416, clk, rst, out_s417, out_e417, result417);
PE P418(out_s354, out_e417, clk, rst, out_s418, out_e418, result418);
PE P419(out_s355, out_e418, clk, rst, out_s419, out_e419, result419);
PE P420(out_s356, out_e419, clk, rst, out_s420, out_e420, result420);
PE P421(out_s357, out_e420, clk, rst, out_s421, out_e421, result421);
PE P422(out_s358, out_e421, clk, rst, out_s422, out_e422, result422);
PE P423(out_s359, out_e422, clk, rst, out_s423, out_e423, result423);
PE P424(out_s360, out_e423, clk, rst, out_s424, out_e424, result424);
PE P425(out_s361, out_e424, clk, rst, out_s425, out_e425, result425);
PE P426(out_s362, out_e425, clk, rst, out_s426, out_e426, result426);
PE P427(out_s363, out_e426, clk, rst, out_s427, out_e427, result427);
PE P428(out_s364, out_e427, clk, rst, out_s428, out_e428, result428);
PE P429(out_s365, out_e428, clk, rst, out_s429, out_e429, result429);
PE P430(out_s366, out_e429, clk, rst, out_s430, out_e430, result430);
PE P431(out_s367, out_e430, clk, rst, out_s431, out_e431, result431);
PE P432(out_s368, out_e431, clk, rst, out_s432, out_e432, result432);
PE P433(out_s369, out_e432, clk, rst, out_s433, out_e433, result433);
PE P434(out_s370, out_e433, clk, rst, out_s434, out_e434, result434);
PE P435(out_s371, out_e434, clk, rst, out_s435, out_e435, result435);
PE P436(out_s372, out_e435, clk, rst, out_s436, out_e436, result436);
PE P437(out_s373, out_e436, clk, rst, out_s437, out_e437, result437);
PE P438(out_s374, out_e437, clk, rst, out_s438, out_e438, result438);
PE P439(out_s375, out_e438, clk, rst, out_s439, out_e439, result439);
PE P440(out_s376, out_e439, clk, rst, out_s440, out_e440, result440);
PE P441(out_s377, out_e440, clk, rst, out_s441, out_e441, result441);
PE P442(out_s378, out_e441, clk, rst, out_s442, out_e442, result442);
PE P443(out_s379, out_e442, clk, rst, out_s443, out_e443, result443);
PE P444(out_s380, out_e443, clk, rst, out_s444, out_e444, result444);
PE P445(out_s381, out_e444, clk, rst, out_s445, out_e445, result445);
PE P446(out_s382, out_e445, clk, rst, out_s446, out_e446, result446);
PE P447(out_s383, out_e446, clk, rst, out_s447, out_e447, result447);

PE P449(out_s385, out_e448, clk, rst, out_s449, out_e449, result449);
PE P450(out_s386, out_e449, clk, rst, out_s450, out_e450, result450);
PE P451(out_s387, out_e450, clk, rst, out_s451, out_e451, result451);
PE P452(out_s388, out_e451, clk, rst, out_s452, out_e452, result452);
PE P453(out_s389, out_e452, clk, rst, out_s453, out_e453, result453);
PE P454(out_s390, out_e453, clk, rst, out_s454, out_e454, result454);
PE P455(out_s391, out_e454, clk, rst, out_s455, out_e455, result455);
PE P456(out_s392, out_e455, clk, rst, out_s456, out_e456, result456);
PE P457(out_s393, out_e456, clk, rst, out_s457, out_e457, result457);
PE P458(out_s394, out_e457, clk, rst, out_s458, out_e458, result458);
PE P459(out_s395, out_e458, clk, rst, out_s459, out_e459, result459);
PE P460(out_s396, out_e459, clk, rst, out_s460, out_e460, result460);
PE P461(out_s397, out_e460, clk, rst, out_s461, out_e461, result461);
PE P462(out_s398, out_e461, clk, rst, out_s462, out_e462, result462);
PE P463(out_s399, out_e462, clk, rst, out_s463, out_e463, result463);
PE P464(out_s400, out_e463, clk, rst, out_s464, out_e464, result464);
PE P465(out_s401, out_e464, clk, rst, out_s465, out_e465, result465);
PE P466(out_s402, out_e465, clk, rst, out_s466, out_e466, result466);
PE P467(out_s403, out_e466, clk, rst, out_s467, out_e467, result467);
PE P468(out_s404, out_e467, clk, rst, out_s468, out_e468, result468);
PE P469(out_s405, out_e468, clk, rst, out_s469, out_e469, result469);
PE P470(out_s406, out_e469, clk, rst, out_s470, out_e470, result470);
PE P471(out_s407, out_e470, clk, rst, out_s471, out_e471, result471);
PE P472(out_s408, out_e471, clk, rst, out_s472, out_e472, result472);
PE P473(out_s409, out_e472, clk, rst, out_s473, out_e473, result473);
PE P474(out_s410, out_e473, clk, rst, out_s474, out_e474, result474);
PE P475(out_s411, out_e474, clk, rst, out_s475, out_e475, result475);
PE P476(out_s412, out_e475, clk, rst, out_s476, out_e476, result476);
PE P477(out_s413, out_e476, clk, rst, out_s477, out_e477, result477);
PE P478(out_s414, out_e477, clk, rst, out_s478, out_e478, result478);
PE P479(out_s415, out_e478, clk, rst, out_s479, out_e479, result479);
PE P480(out_s416, out_e479, clk, rst, out_s480, out_e480, result480);
PE P481(out_s417, out_e480, clk, rst, out_s481, out_e481, result481);
PE P482(out_s418, out_e481, clk, rst, out_s482, out_e482, result482);
PE P483(out_s419, out_e482, clk, rst, out_s483, out_e483, result483);
PE P484(out_s420, out_e483, clk, rst, out_s484, out_e484, result484);
PE P485(out_s421, out_e484, clk, rst, out_s485, out_e485, result485);
PE P486(out_s422, out_e485, clk, rst, out_s486, out_e486, result486);
PE P487(out_s423, out_e486, clk, rst, out_s487, out_e487, result487);
PE P488(out_s424, out_e487, clk, rst, out_s488, out_e488, result488);
PE P489(out_s425, out_e488, clk, rst, out_s489, out_e489, result489);
PE P490(out_s426, out_e489, clk, rst, out_s490, out_e490, result490);
PE P491(out_s427, out_e490, clk, rst, out_s491, out_e491, result491);
PE P492(out_s428, out_e491, clk, rst, out_s492, out_e492, result492);
PE P493(out_s429, out_e492, clk, rst, out_s493, out_e493, result493);
PE P494(out_s430, out_e493, clk, rst, out_s494, out_e494, result494);
PE P495(out_s431, out_e494, clk, rst, out_s495, out_e495, result495);
PE P496(out_s432, out_e495, clk, rst, out_s496, out_e496, result496);
PE P497(out_s433, out_e496, clk, rst, out_s497, out_e497, result497);
PE P498(out_s434, out_e497, clk, rst, out_s498, out_e498, result498);
PE P499(out_s435, out_e498, clk, rst, out_s499, out_e499, result499);
PE P500(out_s436, out_e499, clk, rst, out_s500, out_e500, result500);
PE P501(out_s437, out_e500, clk, rst, out_s501, out_e501, result501);
PE P502(out_s438, out_e501, clk, rst, out_s502, out_e502, result502);
PE P503(out_s439, out_e502, clk, rst, out_s503, out_e503, result503);
PE P504(out_s440, out_e503, clk, rst, out_s504, out_e504, result504);
PE P505(out_s441, out_e504, clk, rst, out_s505, out_e505, result505);
PE P506(out_s442, out_e505, clk, rst, out_s506, out_e506, result506);
PE P507(out_s443, out_e506, clk, rst, out_s507, out_e507, result507);
PE P508(out_s444, out_e507, clk, rst, out_s508, out_e508, result508);
PE P509(out_s445, out_e508, clk, rst, out_s509, out_e509, result509);
PE P510(out_s446, out_e509, clk, rst, out_s510, out_e510, result510);
PE P511(out_s447, out_e510, clk, rst, out_s511, out_e511, result511);

PE P513(out_s449, out_e512, clk, rst, out_s513, out_e513, result513);
PE P514(out_s450, out_e513, clk, rst, out_s514, out_e514, result514);
PE P515(out_s451, out_e514, clk, rst, out_s515, out_e515, result515);
PE P516(out_s452, out_e515, clk, rst, out_s516, out_e516, result516);
PE P517(out_s453, out_e516, clk, rst, out_s517, out_e517, result517);
PE P518(out_s454, out_e517, clk, rst, out_s518, out_e518, result518);
PE P519(out_s455, out_e518, clk, rst, out_s519, out_e519, result519);
PE P520(out_s456, out_e519, clk, rst, out_s520, out_e520, result520);
PE P521(out_s457, out_e520, clk, rst, out_s521, out_e521, result521);
PE P522(out_s458, out_e521, clk, rst, out_s522, out_e522, result522);
PE P523(out_s459, out_e522, clk, rst, out_s523, out_e523, result523);
PE P524(out_s460, out_e523, clk, rst, out_s524, out_e524, result524);
PE P525(out_s461, out_e524, clk, rst, out_s525, out_e525, result525);
PE P526(out_s462, out_e525, clk, rst, out_s526, out_e526, result526);
PE P527(out_s463, out_e526, clk, rst, out_s527, out_e527, result527);
PE P528(out_s464, out_e527, clk, rst, out_s528, out_e528, result528);
PE P529(out_s465, out_e528, clk, rst, out_s529, out_e529, result529);
PE P530(out_s466, out_e529, clk, rst, out_s530, out_e530, result530);
PE P531(out_s467, out_e530, clk, rst, out_s531, out_e531, result531);
PE P532(out_s468, out_e531, clk, rst, out_s532, out_e532, result532);
PE P533(out_s469, out_e532, clk, rst, out_s533, out_e533, result533);
PE P534(out_s470, out_e533, clk, rst, out_s534, out_e534, result534);
PE P535(out_s471, out_e534, clk, rst, out_s535, out_e535, result535);
PE P536(out_s472, out_e535, clk, rst, out_s536, out_e536, result536);
PE P537(out_s473, out_e536, clk, rst, out_s537, out_e537, result537);
PE P538(out_s474, out_e537, clk, rst, out_s538, out_e538, result538);
PE P539(out_s475, out_e538, clk, rst, out_s539, out_e539, result539);
PE P540(out_s476, out_e539, clk, rst, out_s540, out_e540, result540);
PE P541(out_s477, out_e540, clk, rst, out_s541, out_e541, result541);
PE P542(out_s478, out_e541, clk, rst, out_s542, out_e542, result542);
PE P543(out_s479, out_e542, clk, rst, out_s543, out_e543, result543);
PE P544(out_s480, out_e543, clk, rst, out_s544, out_e544, result544);
PE P545(out_s481, out_e544, clk, rst, out_s545, out_e545, result545);
PE P546(out_s482, out_e545, clk, rst, out_s546, out_e546, result546);
PE P547(out_s483, out_e546, clk, rst, out_s547, out_e547, result547);
PE P548(out_s484, out_e547, clk, rst, out_s548, out_e548, result548);
PE P549(out_s485, out_e548, clk, rst, out_s549, out_e549, result549);
PE P550(out_s486, out_e549, clk, rst, out_s550, out_e550, result550);
PE P551(out_s487, out_e550, clk, rst, out_s551, out_e551, result551);
PE P552(out_s488, out_e551, clk, rst, out_s552, out_e552, result552);
PE P553(out_s489, out_e552, clk, rst, out_s553, out_e553, result553);
PE P554(out_s490, out_e553, clk, rst, out_s554, out_e554, result554);
PE P555(out_s491, out_e554, clk, rst, out_s555, out_e555, result555);
PE P556(out_s492, out_e555, clk, rst, out_s556, out_e556, result556);
PE P557(out_s493, out_e556, clk, rst, out_s557, out_e557, result557);
PE P558(out_s494, out_e557, clk, rst, out_s558, out_e558, result558);
PE P559(out_s495, out_e558, clk, rst, out_s559, out_e559, result559);
PE P560(out_s496, out_e559, clk, rst, out_s560, out_e560, result560);
PE P561(out_s497, out_e560, clk, rst, out_s561, out_e561, result561);
PE P562(out_s498, out_e561, clk, rst, out_s562, out_e562, result562);
PE P563(out_s499, out_e562, clk, rst, out_s563, out_e563, result563);
PE P564(out_s500, out_e563, clk, rst, out_s564, out_e564, result564);
PE P565(out_s501, out_e564, clk, rst, out_s565, out_e565, result565);
PE P566(out_s502, out_e565, clk, rst, out_s566, out_e566, result566);
PE P567(out_s503, out_e566, clk, rst, out_s567, out_e567, result567);
PE P568(out_s504, out_e567, clk, rst, out_s568, out_e568, result568);
PE P569(out_s505, out_e568, clk, rst, out_s569, out_e569, result569);
PE P570(out_s506, out_e569, clk, rst, out_s570, out_e570, result570);
PE P571(out_s507, out_e570, clk, rst, out_s571, out_e571, result571);
PE P572(out_s508, out_e571, clk, rst, out_s572, out_e572, result572);
PE P573(out_s509, out_e572, clk, rst, out_s573, out_e573, result573);
PE P574(out_s510, out_e573, clk, rst, out_s574, out_e574, result574);
PE P575(out_s511, out_e574, clk, rst, out_s575, out_e575, result575);

PE P577(out_s513, out_e576, clk, rst, out_s577, out_e577, result577);
PE P578(out_s514, out_e577, clk, rst, out_s578, out_e578, result578);
PE P579(out_s515, out_e578, clk, rst, out_s579, out_e579, result579);
PE P580(out_s516, out_e579, clk, rst, out_s580, out_e580, result580);
PE P581(out_s517, out_e580, clk, rst, out_s581, out_e581, result581);
PE P582(out_s518, out_e581, clk, rst, out_s582, out_e582, result582);
PE P583(out_s519, out_e582, clk, rst, out_s583, out_e583, result583);
PE P584(out_s520, out_e583, clk, rst, out_s584, out_e584, result584);
PE P585(out_s521, out_e584, clk, rst, out_s585, out_e585, result585);
PE P586(out_s522, out_e585, clk, rst, out_s586, out_e586, result586);
PE P587(out_s523, out_e586, clk, rst, out_s587, out_e587, result587);
PE P588(out_s524, out_e587, clk, rst, out_s588, out_e588, result588);
PE P589(out_s525, out_e588, clk, rst, out_s589, out_e589, result589);
PE P590(out_s526, out_e589, clk, rst, out_s590, out_e590, result590);
PE P591(out_s527, out_e590, clk, rst, out_s591, out_e591, result591);
PE P592(out_s528, out_e591, clk, rst, out_s592, out_e592, result592);
PE P593(out_s529, out_e592, clk, rst, out_s593, out_e593, result593);
PE P594(out_s530, out_e593, clk, rst, out_s594, out_e594, result594);
PE P595(out_s531, out_e594, clk, rst, out_s595, out_e595, result595);
PE P596(out_s532, out_e595, clk, rst, out_s596, out_e596, result596);
PE P597(out_s533, out_e596, clk, rst, out_s597, out_e597, result597);
PE P598(out_s534, out_e597, clk, rst, out_s598, out_e598, result598);
PE P599(out_s535, out_e598, clk, rst, out_s599, out_e599, result599);
PE P600(out_s536, out_e599, clk, rst, out_s600, out_e600, result600);
PE P601(out_s537, out_e600, clk, rst, out_s601, out_e601, result601);
PE P602(out_s538, out_e601, clk, rst, out_s602, out_e602, result602);
PE P603(out_s539, out_e602, clk, rst, out_s603, out_e603, result603);
PE P604(out_s540, out_e603, clk, rst, out_s604, out_e604, result604);
PE P605(out_s541, out_e604, clk, rst, out_s605, out_e605, result605);
PE P606(out_s542, out_e605, clk, rst, out_s606, out_e606, result606);
PE P607(out_s543, out_e606, clk, rst, out_s607, out_e607, result607);
PE P608(out_s544, out_e607, clk, rst, out_s608, out_e608, result608);
PE P609(out_s545, out_e608, clk, rst, out_s609, out_e609, result609);
PE P610(out_s546, out_e609, clk, rst, out_s610, out_e610, result610);
PE P611(out_s547, out_e610, clk, rst, out_s611, out_e611, result611);
PE P612(out_s548, out_e611, clk, rst, out_s612, out_e612, result612);
PE P613(out_s549, out_e612, clk, rst, out_s613, out_e613, result613);
PE P614(out_s550, out_e613, clk, rst, out_s614, out_e614, result614);
PE P615(out_s551, out_e614, clk, rst, out_s615, out_e615, result615);
PE P616(out_s552, out_e615, clk, rst, out_s616, out_e616, result616);
PE P617(out_s553, out_e616, clk, rst, out_s617, out_e617, result617);
PE P618(out_s554, out_e617, clk, rst, out_s618, out_e618, result618);
PE P619(out_s555, out_e618, clk, rst, out_s619, out_e619, result619);
PE P620(out_s556, out_e619, clk, rst, out_s620, out_e620, result620);
PE P621(out_s557, out_e620, clk, rst, out_s621, out_e621, result621);
PE P622(out_s558, out_e621, clk, rst, out_s622, out_e622, result622);
PE P623(out_s559, out_e622, clk, rst, out_s623, out_e623, result623);
PE P624(out_s560, out_e623, clk, rst, out_s624, out_e624, result624);
PE P625(out_s561, out_e624, clk, rst, out_s625, out_e625, result625);
PE P626(out_s562, out_e625, clk, rst, out_s626, out_e626, result626);
PE P627(out_s563, out_e626, clk, rst, out_s627, out_e627, result627);
PE P628(out_s564, out_e627, clk, rst, out_s628, out_e628, result628);
PE P629(out_s565, out_e628, clk, rst, out_s629, out_e629, result629);
PE P630(out_s566, out_e629, clk, rst, out_s630, out_e630, result630);
PE P631(out_s567, out_e630, clk, rst, out_s631, out_e631, result631);
PE P632(out_s568, out_e631, clk, rst, out_s632, out_e632, result632);
PE P633(out_s569, out_e632, clk, rst, out_s633, out_e633, result633);
PE P634(out_s570, out_e633, clk, rst, out_s634, out_e634, result634);
PE P635(out_s571, out_e634, clk, rst, out_s635, out_e635, result635);
PE P636(out_s572, out_e635, clk, rst, out_s636, out_e636, result636);
PE P637(out_s573, out_e636, clk, rst, out_s637, out_e637, result637);
PE P638(out_s574, out_e637, clk, rst, out_s638, out_e638, result638);
PE P639(out_s575, out_e638, clk, rst, out_s639, out_e639, result639);

PE P641(out_s577, out_e640, clk, rst, out_s641, out_e641, result641);
PE P642(out_s578, out_e641, clk, rst, out_s642, out_e642, result642);
PE P643(out_s579, out_e642, clk, rst, out_s643, out_e643, result643);
PE P644(out_s580, out_e643, clk, rst, out_s644, out_e644, result644);
PE P645(out_s581, out_e644, clk, rst, out_s645, out_e645, result645);
PE P646(out_s582, out_e645, clk, rst, out_s646, out_e646, result646);
PE P647(out_s583, out_e646, clk, rst, out_s647, out_e647, result647);
PE P648(out_s584, out_e647, clk, rst, out_s648, out_e648, result648);
PE P649(out_s585, out_e648, clk, rst, out_s649, out_e649, result649);
PE P650(out_s586, out_e649, clk, rst, out_s650, out_e650, result650);
PE P651(out_s587, out_e650, clk, rst, out_s651, out_e651, result651);
PE P652(out_s588, out_e651, clk, rst, out_s652, out_e652, result652);
PE P653(out_s589, out_e652, clk, rst, out_s653, out_e653, result653);
PE P654(out_s590, out_e653, clk, rst, out_s654, out_e654, result654);
PE P655(out_s591, out_e654, clk, rst, out_s655, out_e655, result655);
PE P656(out_s592, out_e655, clk, rst, out_s656, out_e656, result656);
PE P657(out_s593, out_e656, clk, rst, out_s657, out_e657, result657);
PE P658(out_s594, out_e657, clk, rst, out_s658, out_e658, result658);
PE P659(out_s595, out_e658, clk, rst, out_s659, out_e659, result659);
PE P660(out_s596, out_e659, clk, rst, out_s660, out_e660, result660);
PE P661(out_s597, out_e660, clk, rst, out_s661, out_e661, result661);
PE P662(out_s598, out_e661, clk, rst, out_s662, out_e662, result662);
PE P663(out_s599, out_e662, clk, rst, out_s663, out_e663, result663);
PE P664(out_s600, out_e663, clk, rst, out_s664, out_e664, result664);
PE P665(out_s601, out_e664, clk, rst, out_s665, out_e665, result665);
PE P666(out_s602, out_e665, clk, rst, out_s666, out_e666, result666);
PE P667(out_s603, out_e666, clk, rst, out_s667, out_e667, result667);
PE P668(out_s604, out_e667, clk, rst, out_s668, out_e668, result668);
PE P669(out_s605, out_e668, clk, rst, out_s669, out_e669, result669);
PE P670(out_s606, out_e669, clk, rst, out_s670, out_e670, result670);
PE P671(out_s607, out_e670, clk, rst, out_s671, out_e671, result671);
PE P672(out_s608, out_e671, clk, rst, out_s672, out_e672, result672);
PE P673(out_s609, out_e672, clk, rst, out_s673, out_e673, result673);
PE P674(out_s610, out_e673, clk, rst, out_s674, out_e674, result674);
PE P675(out_s611, out_e674, clk, rst, out_s675, out_e675, result675);
PE P676(out_s612, out_e675, clk, rst, out_s676, out_e676, result676);
PE P677(out_s613, out_e676, clk, rst, out_s677, out_e677, result677);
PE P678(out_s614, out_e677, clk, rst, out_s678, out_e678, result678);
PE P679(out_s615, out_e678, clk, rst, out_s679, out_e679, result679);
PE P680(out_s616, out_e679, clk, rst, out_s680, out_e680, result680);
PE P681(out_s617, out_e680, clk, rst, out_s681, out_e681, result681);
PE P682(out_s618, out_e681, clk, rst, out_s682, out_e682, result682);
PE P683(out_s619, out_e682, clk, rst, out_s683, out_e683, result683);
PE P684(out_s620, out_e683, clk, rst, out_s684, out_e684, result684);
PE P685(out_s621, out_e684, clk, rst, out_s685, out_e685, result685);
PE P686(out_s622, out_e685, clk, rst, out_s686, out_e686, result686);
PE P687(out_s623, out_e686, clk, rst, out_s687, out_e687, result687);
PE P688(out_s624, out_e687, clk, rst, out_s688, out_e688, result688);
PE P689(out_s625, out_e688, clk, rst, out_s689, out_e689, result689);
PE P690(out_s626, out_e689, clk, rst, out_s690, out_e690, result690);
PE P691(out_s627, out_e690, clk, rst, out_s691, out_e691, result691);
PE P692(out_s628, out_e691, clk, rst, out_s692, out_e692, result692);
PE P693(out_s629, out_e692, clk, rst, out_s693, out_e693, result693);
PE P694(out_s630, out_e693, clk, rst, out_s694, out_e694, result694);
PE P695(out_s631, out_e694, clk, rst, out_s695, out_e695, result695);
PE P696(out_s632, out_e695, clk, rst, out_s696, out_e696, result696);
PE P697(out_s633, out_e696, clk, rst, out_s697, out_e697, result697);
PE P698(out_s634, out_e697, clk, rst, out_s698, out_e698, result698);
PE P699(out_s635, out_e698, clk, rst, out_s699, out_e699, result699);
PE P700(out_s636, out_e699, clk, rst, out_s700, out_e700, result700);
PE P701(out_s637, out_e700, clk, rst, out_s701, out_e701, result701);
PE P702(out_s638, out_e701, clk, rst, out_s702, out_e702, result702);
PE P703(out_s639, out_e702, clk, rst, out_s703, out_e703, result703);

PE P705(out_s641, out_e704, clk, rst, out_s705, out_e705, result705);
PE P706(out_s642, out_e705, clk, rst, out_s706, out_e706, result706);
PE P707(out_s643, out_e706, clk, rst, out_s707, out_e707, result707);
PE P708(out_s644, out_e707, clk, rst, out_s708, out_e708, result708);
PE P709(out_s645, out_e708, clk, rst, out_s709, out_e709, result709);
PE P710(out_s646, out_e709, clk, rst, out_s710, out_e710, result710);
PE P711(out_s647, out_e710, clk, rst, out_s711, out_e711, result711);
PE P712(out_s648, out_e711, clk, rst, out_s712, out_e712, result712);
PE P713(out_s649, out_e712, clk, rst, out_s713, out_e713, result713);
PE P714(out_s650, out_e713, clk, rst, out_s714, out_e714, result714);
PE P715(out_s651, out_e714, clk, rst, out_s715, out_e715, result715);
PE P716(out_s652, out_e715, clk, rst, out_s716, out_e716, result716);
PE P717(out_s653, out_e716, clk, rst, out_s717, out_e717, result717);
PE P718(out_s654, out_e717, clk, rst, out_s718, out_e718, result718);
PE P719(out_s655, out_e718, clk, rst, out_s719, out_e719, result719);
PE P720(out_s656, out_e719, clk, rst, out_s720, out_e720, result720);
PE P721(out_s657, out_e720, clk, rst, out_s721, out_e721, result721);
PE P722(out_s658, out_e721, clk, rst, out_s722, out_e722, result722);
PE P723(out_s659, out_e722, clk, rst, out_s723, out_e723, result723);
PE P724(out_s660, out_e723, clk, rst, out_s724, out_e724, result724);
PE P725(out_s661, out_e724, clk, rst, out_s725, out_e725, result725);
PE P726(out_s662, out_e725, clk, rst, out_s726, out_e726, result726);
PE P727(out_s663, out_e726, clk, rst, out_s727, out_e727, result727);
PE P728(out_s664, out_e727, clk, rst, out_s728, out_e728, result728);
PE P729(out_s665, out_e728, clk, rst, out_s729, out_e729, result729);
PE P730(out_s666, out_e729, clk, rst, out_s730, out_e730, result730);
PE P731(out_s667, out_e730, clk, rst, out_s731, out_e731, result731);
PE P732(out_s668, out_e731, clk, rst, out_s732, out_e732, result732);
PE P733(out_s669, out_e732, clk, rst, out_s733, out_e733, result733);
PE P734(out_s670, out_e733, clk, rst, out_s734, out_e734, result734);
PE P735(out_s671, out_e734, clk, rst, out_s735, out_e735, result735);
PE P736(out_s672, out_e735, clk, rst, out_s736, out_e736, result736);
PE P737(out_s673, out_e736, clk, rst, out_s737, out_e737, result737);
PE P738(out_s674, out_e737, clk, rst, out_s738, out_e738, result738);
PE P739(out_s675, out_e738, clk, rst, out_s739, out_e739, result739);
PE P740(out_s676, out_e739, clk, rst, out_s740, out_e740, result740);
PE P741(out_s677, out_e740, clk, rst, out_s741, out_e741, result741);
PE P742(out_s678, out_e741, clk, rst, out_s742, out_e742, result742);
PE P743(out_s679, out_e742, clk, rst, out_s743, out_e743, result743);
PE P744(out_s680, out_e743, clk, rst, out_s744, out_e744, result744);
PE P745(out_s681, out_e744, clk, rst, out_s745, out_e745, result745);
PE P746(out_s682, out_e745, clk, rst, out_s746, out_e746, result746);
PE P747(out_s683, out_e746, clk, rst, out_s747, out_e747, result747);
PE P748(out_s684, out_e747, clk, rst, out_s748, out_e748, result748);
PE P749(out_s685, out_e748, clk, rst, out_s749, out_e749, result749);
PE P750(out_s686, out_e749, clk, rst, out_s750, out_e750, result750);
PE P751(out_s687, out_e750, clk, rst, out_s751, out_e751, result751);
PE P752(out_s688, out_e751, clk, rst, out_s752, out_e752, result752);
PE P753(out_s689, out_e752, clk, rst, out_s753, out_e753, result753);
PE P754(out_s690, out_e753, clk, rst, out_s754, out_e754, result754);
PE P755(out_s691, out_e754, clk, rst, out_s755, out_e755, result755);
PE P756(out_s692, out_e755, clk, rst, out_s756, out_e756, result756);
PE P757(out_s693, out_e756, clk, rst, out_s757, out_e757, result757);
PE P758(out_s694, out_e757, clk, rst, out_s758, out_e758, result758);
PE P759(out_s695, out_e758, clk, rst, out_s759, out_e759, result759);
PE P760(out_s696, out_e759, clk, rst, out_s760, out_e760, result760);
PE P761(out_s697, out_e760, clk, rst, out_s761, out_e761, result761);
PE P762(out_s698, out_e761, clk, rst, out_s762, out_e762, result762);
PE P763(out_s699, out_e762, clk, rst, out_s763, out_e763, result763);
PE P764(out_s700, out_e763, clk, rst, out_s764, out_e764, result764);
PE P765(out_s701, out_e764, clk, rst, out_s765, out_e765, result765);
PE P766(out_s702, out_e765, clk, rst, out_s766, out_e766, result766);
PE P767(out_s703, out_e766, clk, rst, out_s767, out_e767, result767);

PE P769(out_s705, out_e768, clk, rst, out_s769, out_e769, result769);
PE P770(out_s706, out_e769, clk, rst, out_s770, out_e770, result770);
PE P771(out_s707, out_e770, clk, rst, out_s771, out_e771, result771);
PE P772(out_s708, out_e771, clk, rst, out_s772, out_e772, result772);
PE P773(out_s709, out_e772, clk, rst, out_s773, out_e773, result773);
PE P774(out_s710, out_e773, clk, rst, out_s774, out_e774, result774);
PE P775(out_s711, out_e774, clk, rst, out_s775, out_e775, result775);
PE P776(out_s712, out_e775, clk, rst, out_s776, out_e776, result776);
PE P777(out_s713, out_e776, clk, rst, out_s777, out_e777, result777);
PE P778(out_s714, out_e777, clk, rst, out_s778, out_e778, result778);
PE P779(out_s715, out_e778, clk, rst, out_s779, out_e779, result779);
PE P780(out_s716, out_e779, clk, rst, out_s780, out_e780, result780);
PE P781(out_s717, out_e780, clk, rst, out_s781, out_e781, result781);
PE P782(out_s718, out_e781, clk, rst, out_s782, out_e782, result782);
PE P783(out_s719, out_e782, clk, rst, out_s783, out_e783, result783);
PE P784(out_s720, out_e783, clk, rst, out_s784, out_e784, result784);
PE P785(out_s721, out_e784, clk, rst, out_s785, out_e785, result785);
PE P786(out_s722, out_e785, clk, rst, out_s786, out_e786, result786);
PE P787(out_s723, out_e786, clk, rst, out_s787, out_e787, result787);
PE P788(out_s724, out_e787, clk, rst, out_s788, out_e788, result788);
PE P789(out_s725, out_e788, clk, rst, out_s789, out_e789, result789);
PE P790(out_s726, out_e789, clk, rst, out_s790, out_e790, result790);
PE P791(out_s727, out_e790, clk, rst, out_s791, out_e791, result791);
PE P792(out_s728, out_e791, clk, rst, out_s792, out_e792, result792);
PE P793(out_s729, out_e792, clk, rst, out_s793, out_e793, result793);
PE P794(out_s730, out_e793, clk, rst, out_s794, out_e794, result794);
PE P795(out_s731, out_e794, clk, rst, out_s795, out_e795, result795);
PE P796(out_s732, out_e795, clk, rst, out_s796, out_e796, result796);
PE P797(out_s733, out_e796, clk, rst, out_s797, out_e797, result797);
PE P798(out_s734, out_e797, clk, rst, out_s798, out_e798, result798);
PE P799(out_s735, out_e798, clk, rst, out_s799, out_e799, result799);
PE P800(out_s736, out_e799, clk, rst, out_s800, out_e800, result800);
PE P801(out_s737, out_e800, clk, rst, out_s801, out_e801, result801);
PE P802(out_s738, out_e801, clk, rst, out_s802, out_e802, result802);
PE P803(out_s739, out_e802, clk, rst, out_s803, out_e803, result803);
PE P804(out_s740, out_e803, clk, rst, out_s804, out_e804, result804);
PE P805(out_s741, out_e804, clk, rst, out_s805, out_e805, result805);
PE P806(out_s742, out_e805, clk, rst, out_s806, out_e806, result806);
PE P807(out_s743, out_e806, clk, rst, out_s807, out_e807, result807);
PE P808(out_s744, out_e807, clk, rst, out_s808, out_e808, result808);
PE P809(out_s745, out_e808, clk, rst, out_s809, out_e809, result809);
PE P810(out_s746, out_e809, clk, rst, out_s810, out_e810, result810);
PE P811(out_s747, out_e810, clk, rst, out_s811, out_e811, result811);
PE P812(out_s748, out_e811, clk, rst, out_s812, out_e812, result812);
PE P813(out_s749, out_e812, clk, rst, out_s813, out_e813, result813);
PE P814(out_s750, out_e813, clk, rst, out_s814, out_e814, result814);
PE P815(out_s751, out_e814, clk, rst, out_s815, out_e815, result815);
PE P816(out_s752, out_e815, clk, rst, out_s816, out_e816, result816);
PE P817(out_s753, out_e816, clk, rst, out_s817, out_e817, result817);
PE P818(out_s754, out_e817, clk, rst, out_s818, out_e818, result818);
PE P819(out_s755, out_e818, clk, rst, out_s819, out_e819, result819);
PE P820(out_s756, out_e819, clk, rst, out_s820, out_e820, result820);
PE P821(out_s757, out_e820, clk, rst, out_s821, out_e821, result821);
PE P822(out_s758, out_e821, clk, rst, out_s822, out_e822, result822);
PE P823(out_s759, out_e822, clk, rst, out_s823, out_e823, result823);
PE P824(out_s760, out_e823, clk, rst, out_s824, out_e824, result824);
PE P825(out_s761, out_e824, clk, rst, out_s825, out_e825, result825);
PE P826(out_s762, out_e825, clk, rst, out_s826, out_e826, result826);
PE P827(out_s763, out_e826, clk, rst, out_s827, out_e827, result827);
PE P828(out_s764, out_e827, clk, rst, out_s828, out_e828, result828);
PE P829(out_s765, out_e828, clk, rst, out_s829, out_e829, result829);
PE P830(out_s766, out_e829, clk, rst, out_s830, out_e830, result830);
PE P831(out_s767, out_e830, clk, rst, out_s831, out_e831, result831);

PE P833(out_s769, out_e832, clk, rst, out_s833, out_e833, result833);
PE P834(out_s770, out_e833, clk, rst, out_s834, out_e834, result834);
PE P835(out_s771, out_e834, clk, rst, out_s835, out_e835, result835);
PE P836(out_s772, out_e835, clk, rst, out_s836, out_e836, result836);
PE P837(out_s773, out_e836, clk, rst, out_s837, out_e837, result837);
PE P838(out_s774, out_e837, clk, rst, out_s838, out_e838, result838);
PE P839(out_s775, out_e838, clk, rst, out_s839, out_e839, result839);
PE P840(out_s776, out_e839, clk, rst, out_s840, out_e840, result840);
PE P841(out_s777, out_e840, clk, rst, out_s841, out_e841, result841);
PE P842(out_s778, out_e841, clk, rst, out_s842, out_e842, result842);
PE P843(out_s779, out_e842, clk, rst, out_s843, out_e843, result843);
PE P844(out_s780, out_e843, clk, rst, out_s844, out_e844, result844);
PE P845(out_s781, out_e844, clk, rst, out_s845, out_e845, result845);
PE P846(out_s782, out_e845, clk, rst, out_s846, out_e846, result846);
PE P847(out_s783, out_e846, clk, rst, out_s847, out_e847, result847);
PE P848(out_s784, out_e847, clk, rst, out_s848, out_e848, result848);
PE P849(out_s785, out_e848, clk, rst, out_s849, out_e849, result849);
PE P850(out_s786, out_e849, clk, rst, out_s850, out_e850, result850);
PE P851(out_s787, out_e850, clk, rst, out_s851, out_e851, result851);
PE P852(out_s788, out_e851, clk, rst, out_s852, out_e852, result852);
PE P853(out_s789, out_e852, clk, rst, out_s853, out_e853, result853);
PE P854(out_s790, out_e853, clk, rst, out_s854, out_e854, result854);
PE P855(out_s791, out_e854, clk, rst, out_s855, out_e855, result855);
PE P856(out_s792, out_e855, clk, rst, out_s856, out_e856, result856);
PE P857(out_s793, out_e856, clk, rst, out_s857, out_e857, result857);
PE P858(out_s794, out_e857, clk, rst, out_s858, out_e858, result858);
PE P859(out_s795, out_e858, clk, rst, out_s859, out_e859, result859);
PE P860(out_s796, out_e859, clk, rst, out_s860, out_e860, result860);
PE P861(out_s797, out_e860, clk, rst, out_s861, out_e861, result861);
PE P862(out_s798, out_e861, clk, rst, out_s862, out_e862, result862);
PE P863(out_s799, out_e862, clk, rst, out_s863, out_e863, result863);
PE P864(out_s800, out_e863, clk, rst, out_s864, out_e864, result864);
PE P865(out_s801, out_e864, clk, rst, out_s865, out_e865, result865);
PE P866(out_s802, out_e865, clk, rst, out_s866, out_e866, result866);
PE P867(out_s803, out_e866, clk, rst, out_s867, out_e867, result867);
PE P868(out_s804, out_e867, clk, rst, out_s868, out_e868, result868);
PE P869(out_s805, out_e868, clk, rst, out_s869, out_e869, result869);
PE P870(out_s806, out_e869, clk, rst, out_s870, out_e870, result870);
PE P871(out_s807, out_e870, clk, rst, out_s871, out_e871, result871);
PE P872(out_s808, out_e871, clk, rst, out_s872, out_e872, result872);
PE P873(out_s809, out_e872, clk, rst, out_s873, out_e873, result873);
PE P874(out_s810, out_e873, clk, rst, out_s874, out_e874, result874);
PE P875(out_s811, out_e874, clk, rst, out_s875, out_e875, result875);
PE P876(out_s812, out_e875, clk, rst, out_s876, out_e876, result876);
PE P877(out_s813, out_e876, clk, rst, out_s877, out_e877, result877);
PE P878(out_s814, out_e877, clk, rst, out_s878, out_e878, result878);
PE P879(out_s815, out_e878, clk, rst, out_s879, out_e879, result879);
PE P880(out_s816, out_e879, clk, rst, out_s880, out_e880, result880);
PE P881(out_s817, out_e880, clk, rst, out_s881, out_e881, result881);
PE P882(out_s818, out_e881, clk, rst, out_s882, out_e882, result882);
PE P883(out_s819, out_e882, clk, rst, out_s883, out_e883, result883);
PE P884(out_s820, out_e883, clk, rst, out_s884, out_e884, result884);
PE P885(out_s821, out_e884, clk, rst, out_s885, out_e885, result885);
PE P886(out_s822, out_e885, clk, rst, out_s886, out_e886, result886);
PE P887(out_s823, out_e886, clk, rst, out_s887, out_e887, result887);
PE P888(out_s824, out_e887, clk, rst, out_s888, out_e888, result888);
PE P889(out_s825, out_e888, clk, rst, out_s889, out_e889, result889);
PE P890(out_s826, out_e889, clk, rst, out_s890, out_e890, result890);
PE P891(out_s827, out_e890, clk, rst, out_s891, out_e891, result891);
PE P892(out_s828, out_e891, clk, rst, out_s892, out_e892, result892);
PE P893(out_s829, out_e892, clk, rst, out_s893, out_e893, result893);
PE P894(out_s830, out_e893, clk, rst, out_s894, out_e894, result894);
PE P895(out_s831, out_e894, clk, rst, out_s895, out_e895, result895);

PE P897(out_s833, out_e896, clk, rst, out_s897, out_e897, result897);
PE P898(out_s834, out_e897, clk, rst, out_s898, out_e898, result898);
PE P899(out_s835, out_e898, clk, rst, out_s899, out_e899, result899);
PE P900(out_s836, out_e899, clk, rst, out_s900, out_e900, result900);
PE P901(out_s837, out_e900, clk, rst, out_s901, out_e901, result901);
PE P902(out_s838, out_e901, clk, rst, out_s902, out_e902, result902);
PE P903(out_s839, out_e902, clk, rst, out_s903, out_e903, result903);
PE P904(out_s840, out_e903, clk, rst, out_s904, out_e904, result904);
PE P905(out_s841, out_e904, clk, rst, out_s905, out_e905, result905);
PE P906(out_s842, out_e905, clk, rst, out_s906, out_e906, result906);
PE P907(out_s843, out_e906, clk, rst, out_s907, out_e907, result907);
PE P908(out_s844, out_e907, clk, rst, out_s908, out_e908, result908);
PE P909(out_s845, out_e908, clk, rst, out_s909, out_e909, result909);
PE P910(out_s846, out_e909, clk, rst, out_s910, out_e910, result910);
PE P911(out_s847, out_e910, clk, rst, out_s911, out_e911, result911);
PE P912(out_s848, out_e911, clk, rst, out_s912, out_e912, result912);
PE P913(out_s849, out_e912, clk, rst, out_s913, out_e913, result913);
PE P914(out_s850, out_e913, clk, rst, out_s914, out_e914, result914);
PE P915(out_s851, out_e914, clk, rst, out_s915, out_e915, result915);
PE P916(out_s852, out_e915, clk, rst, out_s916, out_e916, result916);
PE P917(out_s853, out_e916, clk, rst, out_s917, out_e917, result917);
PE P918(out_s854, out_e917, clk, rst, out_s918, out_e918, result918);
PE P919(out_s855, out_e918, clk, rst, out_s919, out_e919, result919);
PE P920(out_s856, out_e919, clk, rst, out_s920, out_e920, result920);
PE P921(out_s857, out_e920, clk, rst, out_s921, out_e921, result921);
PE P922(out_s858, out_e921, clk, rst, out_s922, out_e922, result922);
PE P923(out_s859, out_e922, clk, rst, out_s923, out_e923, result923);
PE P924(out_s860, out_e923, clk, rst, out_s924, out_e924, result924);
PE P925(out_s861, out_e924, clk, rst, out_s925, out_e925, result925);
PE P926(out_s862, out_e925, clk, rst, out_s926, out_e926, result926);
PE P927(out_s863, out_e926, clk, rst, out_s927, out_e927, result927);
PE P928(out_s864, out_e927, clk, rst, out_s928, out_e928, result928);
PE P929(out_s865, out_e928, clk, rst, out_s929, out_e929, result929);
PE P930(out_s866, out_e929, clk, rst, out_s930, out_e930, result930);
PE P931(out_s867, out_e930, clk, rst, out_s931, out_e931, result931);
PE P932(out_s868, out_e931, clk, rst, out_s932, out_e932, result932);
PE P933(out_s869, out_e932, clk, rst, out_s933, out_e933, result933);
PE P934(out_s870, out_e933, clk, rst, out_s934, out_e934, result934);
PE P935(out_s871, out_e934, clk, rst, out_s935, out_e935, result935);
PE P936(out_s872, out_e935, clk, rst, out_s936, out_e936, result936);
PE P937(out_s873, out_e936, clk, rst, out_s937, out_e937, result937);
PE P938(out_s874, out_e937, clk, rst, out_s938, out_e938, result938);
PE P939(out_s875, out_e938, clk, rst, out_s939, out_e939, result939);
PE P940(out_s876, out_e939, clk, rst, out_s940, out_e940, result940);
PE P941(out_s877, out_e940, clk, rst, out_s941, out_e941, result941);
PE P942(out_s878, out_e941, clk, rst, out_s942, out_e942, result942);
PE P943(out_s879, out_e942, clk, rst, out_s943, out_e943, result943);
PE P944(out_s880, out_e943, clk, rst, out_s944, out_e944, result944);
PE P945(out_s881, out_e944, clk, rst, out_s945, out_e945, result945);
PE P946(out_s882, out_e945, clk, rst, out_s946, out_e946, result946);
PE P947(out_s883, out_e946, clk, rst, out_s947, out_e947, result947);
PE P948(out_s884, out_e947, clk, rst, out_s948, out_e948, result948);
PE P949(out_s885, out_e948, clk, rst, out_s949, out_e949, result949);
PE P950(out_s886, out_e949, clk, rst, out_s950, out_e950, result950);
PE P951(out_s887, out_e950, clk, rst, out_s951, out_e951, result951);
PE P952(out_s888, out_e951, clk, rst, out_s952, out_e952, result952);
PE P953(out_s889, out_e952, clk, rst, out_s953, out_e953, result953);
PE P954(out_s890, out_e953, clk, rst, out_s954, out_e954, result954);
PE P955(out_s891, out_e954, clk, rst, out_s955, out_e955, result955);
PE P956(out_s892, out_e955, clk, rst, out_s956, out_e956, result956);
PE P957(out_s893, out_e956, clk, rst, out_s957, out_e957, result957);
PE P958(out_s894, out_e957, clk, rst, out_s958, out_e958, result958);
PE P959(out_s895, out_e958, clk, rst, out_s959, out_e959, result959);

PE P961(out_s897, out_e960, clk, rst, out_s961, out_e961, result961);
PE P962(out_s898, out_e961, clk, rst, out_s962, out_e962, result962);
PE P963(out_s899, out_e962, clk, rst, out_s963, out_e963, result963);
PE P964(out_s900, out_e963, clk, rst, out_s964, out_e964, result964);
PE P965(out_s901, out_e964, clk, rst, out_s965, out_e965, result965);
PE P966(out_s902, out_e965, clk, rst, out_s966, out_e966, result966);
PE P967(out_s903, out_e966, clk, rst, out_s967, out_e967, result967);
PE P968(out_s904, out_e967, clk, rst, out_s968, out_e968, result968);
PE P969(out_s905, out_e968, clk, rst, out_s969, out_e969, result969);
PE P970(out_s906, out_e969, clk, rst, out_s970, out_e970, result970);
PE P971(out_s907, out_e970, clk, rst, out_s971, out_e971, result971);
PE P972(out_s908, out_e971, clk, rst, out_s972, out_e972, result972);
PE P973(out_s909, out_e972, clk, rst, out_s973, out_e973, result973);
PE P974(out_s910, out_e973, clk, rst, out_s974, out_e974, result974);
PE P975(out_s911, out_e974, clk, rst, out_s975, out_e975, result975);
PE P976(out_s912, out_e975, clk, rst, out_s976, out_e976, result976);
PE P977(out_s913, out_e976, clk, rst, out_s977, out_e977, result977);
PE P978(out_s914, out_e977, clk, rst, out_s978, out_e978, result978);
PE P979(out_s915, out_e978, clk, rst, out_s979, out_e979, result979);
PE P980(out_s916, out_e979, clk, rst, out_s980, out_e980, result980);
PE P981(out_s917, out_e980, clk, rst, out_s981, out_e981, result981);
PE P982(out_s918, out_e981, clk, rst, out_s982, out_e982, result982);
PE P983(out_s919, out_e982, clk, rst, out_s983, out_e983, result983);
PE P984(out_s920, out_e983, clk, rst, out_s984, out_e984, result984);
PE P985(out_s921, out_e984, clk, rst, out_s985, out_e985, result985);
PE P986(out_s922, out_e985, clk, rst, out_s986, out_e986, result986);
PE P987(out_s923, out_e986, clk, rst, out_s987, out_e987, result987);
PE P988(out_s924, out_e987, clk, rst, out_s988, out_e988, result988);
PE P989(out_s925, out_e988, clk, rst, out_s989, out_e989, result989);
PE P990(out_s926, out_e989, clk, rst, out_s990, out_e990, result990);
PE P991(out_s927, out_e990, clk, rst, out_s991, out_e991, result991);
PE P992(out_s928, out_e991, clk, rst, out_s992, out_e992, result992);
PE P993(out_s929, out_e992, clk, rst, out_s993, out_e993, result993);
PE P994(out_s930, out_e993, clk, rst, out_s994, out_e994, result994);
PE P995(out_s931, out_e994, clk, rst, out_s995, out_e995, result995);
PE P996(out_s932, out_e995, clk, rst, out_s996, out_e996, result996);
PE P997(out_s933, out_e996, clk, rst, out_s997, out_e997, result997);
PE P998(out_s934, out_e997, clk, rst, out_s998, out_e998, result998);
PE P999(out_s935, out_e998, clk, rst, out_s999, out_e999, result999);
PE P1000(out_s936, out_e999, clk, rst, out_s1000, out_e1000, result1000);
PE P1001(out_s937, out_e1000, clk, rst, out_s1001, out_e1001, result1001);
PE P1002(out_s938, out_e1001, clk, rst, out_s1002, out_e1002, result1002);
PE P1003(out_s939, out_e1002, clk, rst, out_s1003, out_e1003, result1003);
PE P1004(out_s940, out_e1003, clk, rst, out_s1004, out_e1004, result1004);
PE P1005(out_s941, out_e1004, clk, rst, out_s1005, out_e1005, result1005);
PE P1006(out_s942, out_e1005, clk, rst, out_s1006, out_e1006, result1006);
PE P1007(out_s943, out_e1006, clk, rst, out_s1007, out_e1007, result1007);
PE P1008(out_s944, out_e1007, clk, rst, out_s1008, out_e1008, result1008);
PE P1009(out_s945, out_e1008, clk, rst, out_s1009, out_e1009, result1009);
PE P1010(out_s946, out_e1009, clk, rst, out_s1010, out_e1010, result1010);
PE P1011(out_s947, out_e1010, clk, rst, out_s1011, out_e1011, result1011);
PE P1012(out_s948, out_e1011, clk, rst, out_s1012, out_e1012, result1012);
PE P1013(out_s949, out_e1012, clk, rst, out_s1013, out_e1013, result1013);
PE P1014(out_s950, out_e1013, clk, rst, out_s1014, out_e1014, result1014);
PE P1015(out_s951, out_e1014, clk, rst, out_s1015, out_e1015, result1015);
PE P1016(out_s952, out_e1015, clk, rst, out_s1016, out_e1016, result1016);
PE P1017(out_s953, out_e1016, clk, rst, out_s1017, out_e1017, result1017);
PE P1018(out_s954, out_e1017, clk, rst, out_s1018, out_e1018, result1018);
PE P1019(out_s955, out_e1018, clk, rst, out_s1019, out_e1019, result1019);
PE P1020(out_s956, out_e1019, clk, rst, out_s1020, out_e1020, result1020);
PE P1021(out_s957, out_e1020, clk, rst, out_s1021, out_e1021, result1021);
PE P1022(out_s958, out_e1021, clk, rst, out_s1022, out_e1022, result1022);
PE P1023(out_s959, out_e1022, clk, rst, out_s1023, out_e1023, result1023);

PE P1025(out_s961, out_e1024, clk, rst, out_s1025, out_e1025, result1025);
PE P1026(out_s962, out_e1025, clk, rst, out_s1026, out_e1026, result1026);
PE P1027(out_s963, out_e1026, clk, rst, out_s1027, out_e1027, result1027);
PE P1028(out_s964, out_e1027, clk, rst, out_s1028, out_e1028, result1028);
PE P1029(out_s965, out_e1028, clk, rst, out_s1029, out_e1029, result1029);
PE P1030(out_s966, out_e1029, clk, rst, out_s1030, out_e1030, result1030);
PE P1031(out_s967, out_e1030, clk, rst, out_s1031, out_e1031, result1031);
PE P1032(out_s968, out_e1031, clk, rst, out_s1032, out_e1032, result1032);
PE P1033(out_s969, out_e1032, clk, rst, out_s1033, out_e1033, result1033);
PE P1034(out_s970, out_e1033, clk, rst, out_s1034, out_e1034, result1034);
PE P1035(out_s971, out_e1034, clk, rst, out_s1035, out_e1035, result1035);
PE P1036(out_s972, out_e1035, clk, rst, out_s1036, out_e1036, result1036);
PE P1037(out_s973, out_e1036, clk, rst, out_s1037, out_e1037, result1037);
PE P1038(out_s974, out_e1037, clk, rst, out_s1038, out_e1038, result1038);
PE P1039(out_s975, out_e1038, clk, rst, out_s1039, out_e1039, result1039);
PE P1040(out_s976, out_e1039, clk, rst, out_s1040, out_e1040, result1040);
PE P1041(out_s977, out_e1040, clk, rst, out_s1041, out_e1041, result1041);
PE P1042(out_s978, out_e1041, clk, rst, out_s1042, out_e1042, result1042);
PE P1043(out_s979, out_e1042, clk, rst, out_s1043, out_e1043, result1043);
PE P1044(out_s980, out_e1043, clk, rst, out_s1044, out_e1044, result1044);
PE P1045(out_s981, out_e1044, clk, rst, out_s1045, out_e1045, result1045);
PE P1046(out_s982, out_e1045, clk, rst, out_s1046, out_e1046, result1046);
PE P1047(out_s983, out_e1046, clk, rst, out_s1047, out_e1047, result1047);
PE P1048(out_s984, out_e1047, clk, rst, out_s1048, out_e1048, result1048);
PE P1049(out_s985, out_e1048, clk, rst, out_s1049, out_e1049, result1049);
PE P1050(out_s986, out_e1049, clk, rst, out_s1050, out_e1050, result1050);
PE P1051(out_s987, out_e1050, clk, rst, out_s1051, out_e1051, result1051);
PE P1052(out_s988, out_e1051, clk, rst, out_s1052, out_e1052, result1052);
PE P1053(out_s989, out_e1052, clk, rst, out_s1053, out_e1053, result1053);
PE P1054(out_s990, out_e1053, clk, rst, out_s1054, out_e1054, result1054);
PE P1055(out_s991, out_e1054, clk, rst, out_s1055, out_e1055, result1055);
PE P1056(out_s992, out_e1055, clk, rst, out_s1056, out_e1056, result1056);
PE P1057(out_s993, out_e1056, clk, rst, out_s1057, out_e1057, result1057);
PE P1058(out_s994, out_e1057, clk, rst, out_s1058, out_e1058, result1058);
PE P1059(out_s995, out_e1058, clk, rst, out_s1059, out_e1059, result1059);
PE P1060(out_s996, out_e1059, clk, rst, out_s1060, out_e1060, result1060);
PE P1061(out_s997, out_e1060, clk, rst, out_s1061, out_e1061, result1061);
PE P1062(out_s998, out_e1061, clk, rst, out_s1062, out_e1062, result1062);
PE P1063(out_s999, out_e1062, clk, rst, out_s1063, out_e1063, result1063);
PE P1064(out_s1000, out_e1063, clk, rst, out_s1064, out_e1064, result1064);
PE P1065(out_s1001, out_e1064, clk, rst, out_s1065, out_e1065, result1065);
PE P1066(out_s1002, out_e1065, clk, rst, out_s1066, out_e1066, result1066);
PE P1067(out_s1003, out_e1066, clk, rst, out_s1067, out_e1067, result1067);
PE P1068(out_s1004, out_e1067, clk, rst, out_s1068, out_e1068, result1068);
PE P1069(out_s1005, out_e1068, clk, rst, out_s1069, out_e1069, result1069);
PE P1070(out_s1006, out_e1069, clk, rst, out_s1070, out_e1070, result1070);
PE P1071(out_s1007, out_e1070, clk, rst, out_s1071, out_e1071, result1071);
PE P1072(out_s1008, out_e1071, clk, rst, out_s1072, out_e1072, result1072);
PE P1073(out_s1009, out_e1072, clk, rst, out_s1073, out_e1073, result1073);
PE P1074(out_s1010, out_e1073, clk, rst, out_s1074, out_e1074, result1074);
PE P1075(out_s1011, out_e1074, clk, rst, out_s1075, out_e1075, result1075);
PE P1076(out_s1012, out_e1075, clk, rst, out_s1076, out_e1076, result1076);
PE P1077(out_s1013, out_e1076, clk, rst, out_s1077, out_e1077, result1077);
PE P1078(out_s1014, out_e1077, clk, rst, out_s1078, out_e1078, result1078);
PE P1079(out_s1015, out_e1078, clk, rst, out_s1079, out_e1079, result1079);
PE P1080(out_s1016, out_e1079, clk, rst, out_s1080, out_e1080, result1080);
PE P1081(out_s1017, out_e1080, clk, rst, out_s1081, out_e1081, result1081);
PE P1082(out_s1018, out_e1081, clk, rst, out_s1082, out_e1082, result1082);
PE P1083(out_s1019, out_e1082, clk, rst, out_s1083, out_e1083, result1083);
PE P1084(out_s1020, out_e1083, clk, rst, out_s1084, out_e1084, result1084);
PE P1085(out_s1021, out_e1084, clk, rst, out_s1085, out_e1085, result1085);
PE P1086(out_s1022, out_e1085, clk, rst, out_s1086, out_e1086, result1086);
PE P1087(out_s1023, out_e1086, clk, rst, out_s1087, out_e1087, result1087);

PE P1089(out_s1025, out_e1088, clk, rst, out_s1089, out_e1089, result1089);
PE P1090(out_s1026, out_e1089, clk, rst, out_s1090, out_e1090, result1090);
PE P1091(out_s1027, out_e1090, clk, rst, out_s1091, out_e1091, result1091);
PE P1092(out_s1028, out_e1091, clk, rst, out_s1092, out_e1092, result1092);
PE P1093(out_s1029, out_e1092, clk, rst, out_s1093, out_e1093, result1093);
PE P1094(out_s1030, out_e1093, clk, rst, out_s1094, out_e1094, result1094);
PE P1095(out_s1031, out_e1094, clk, rst, out_s1095, out_e1095, result1095);
PE P1096(out_s1032, out_e1095, clk, rst, out_s1096, out_e1096, result1096);
PE P1097(out_s1033, out_e1096, clk, rst, out_s1097, out_e1097, result1097);
PE P1098(out_s1034, out_e1097, clk, rst, out_s1098, out_e1098, result1098);
PE P1099(out_s1035, out_e1098, clk, rst, out_s1099, out_e1099, result1099);
PE P1100(out_s1036, out_e1099, clk, rst, out_s1100, out_e1100, result1100);
PE P1101(out_s1037, out_e1100, clk, rst, out_s1101, out_e1101, result1101);
PE P1102(out_s1038, out_e1101, clk, rst, out_s1102, out_e1102, result1102);
PE P1103(out_s1039, out_e1102, clk, rst, out_s1103, out_e1103, result1103);
PE P1104(out_s1040, out_e1103, clk, rst, out_s1104, out_e1104, result1104);
PE P1105(out_s1041, out_e1104, clk, rst, out_s1105, out_e1105, result1105);
PE P1106(out_s1042, out_e1105, clk, rst, out_s1106, out_e1106, result1106);
PE P1107(out_s1043, out_e1106, clk, rst, out_s1107, out_e1107, result1107);
PE P1108(out_s1044, out_e1107, clk, rst, out_s1108, out_e1108, result1108);
PE P1109(out_s1045, out_e1108, clk, rst, out_s1109, out_e1109, result1109);
PE P1110(out_s1046, out_e1109, clk, rst, out_s1110, out_e1110, result1110);
PE P1111(out_s1047, out_e1110, clk, rst, out_s1111, out_e1111, result1111);
PE P1112(out_s1048, out_e1111, clk, rst, out_s1112, out_e1112, result1112);
PE P1113(out_s1049, out_e1112, clk, rst, out_s1113, out_e1113, result1113);
PE P1114(out_s1050, out_e1113, clk, rst, out_s1114, out_e1114, result1114);
PE P1115(out_s1051, out_e1114, clk, rst, out_s1115, out_e1115, result1115);
PE P1116(out_s1052, out_e1115, clk, rst, out_s1116, out_e1116, result1116);
PE P1117(out_s1053, out_e1116, clk, rst, out_s1117, out_e1117, result1117);
PE P1118(out_s1054, out_e1117, clk, rst, out_s1118, out_e1118, result1118);
PE P1119(out_s1055, out_e1118, clk, rst, out_s1119, out_e1119, result1119);
PE P1120(out_s1056, out_e1119, clk, rst, out_s1120, out_e1120, result1120);
PE P1121(out_s1057, out_e1120, clk, rst, out_s1121, out_e1121, result1121);
PE P1122(out_s1058, out_e1121, clk, rst, out_s1122, out_e1122, result1122);
PE P1123(out_s1059, out_e1122, clk, rst, out_s1123, out_e1123, result1123);
PE P1124(out_s1060, out_e1123, clk, rst, out_s1124, out_e1124, result1124);
PE P1125(out_s1061, out_e1124, clk, rst, out_s1125, out_e1125, result1125);
PE P1126(out_s1062, out_e1125, clk, rst, out_s1126, out_e1126, result1126);
PE P1127(out_s1063, out_e1126, clk, rst, out_s1127, out_e1127, result1127);
PE P1128(out_s1064, out_e1127, clk, rst, out_s1128, out_e1128, result1128);
PE P1129(out_s1065, out_e1128, clk, rst, out_s1129, out_e1129, result1129);
PE P1130(out_s1066, out_e1129, clk, rst, out_s1130, out_e1130, result1130);
PE P1131(out_s1067, out_e1130, clk, rst, out_s1131, out_e1131, result1131);
PE P1132(out_s1068, out_e1131, clk, rst, out_s1132, out_e1132, result1132);
PE P1133(out_s1069, out_e1132, clk, rst, out_s1133, out_e1133, result1133);
PE P1134(out_s1070, out_e1133, clk, rst, out_s1134, out_e1134, result1134);
PE P1135(out_s1071, out_e1134, clk, rst, out_s1135, out_e1135, result1135);
PE P1136(out_s1072, out_e1135, clk, rst, out_s1136, out_e1136, result1136);
PE P1137(out_s1073, out_e1136, clk, rst, out_s1137, out_e1137, result1137);
PE P1138(out_s1074, out_e1137, clk, rst, out_s1138, out_e1138, result1138);
PE P1139(out_s1075, out_e1138, clk, rst, out_s1139, out_e1139, result1139);
PE P1140(out_s1076, out_e1139, clk, rst, out_s1140, out_e1140, result1140);
PE P1141(out_s1077, out_e1140, clk, rst, out_s1141, out_e1141, result1141);
PE P1142(out_s1078, out_e1141, clk, rst, out_s1142, out_e1142, result1142);
PE P1143(out_s1079, out_e1142, clk, rst, out_s1143, out_e1143, result1143);
PE P1144(out_s1080, out_e1143, clk, rst, out_s1144, out_e1144, result1144);
PE P1145(out_s1081, out_e1144, clk, rst, out_s1145, out_e1145, result1145);
PE P1146(out_s1082, out_e1145, clk, rst, out_s1146, out_e1146, result1146);
PE P1147(out_s1083, out_e1146, clk, rst, out_s1147, out_e1147, result1147);
PE P1148(out_s1084, out_e1147, clk, rst, out_s1148, out_e1148, result1148);
PE P1149(out_s1085, out_e1148, clk, rst, out_s1149, out_e1149, result1149);
PE P1150(out_s1086, out_e1149, clk, rst, out_s1150, out_e1150, result1150);
PE P1151(out_s1087, out_e1150, clk, rst, out_s1151, out_e1151, result1151);

PE P1153(out_s1089, out_e1152, clk, rst, out_s1153, out_e1153, result1153);
PE P1154(out_s1090, out_e1153, clk, rst, out_s1154, out_e1154, result1154);
PE P1155(out_s1091, out_e1154, clk, rst, out_s1155, out_e1155, result1155);
PE P1156(out_s1092, out_e1155, clk, rst, out_s1156, out_e1156, result1156);
PE P1157(out_s1093, out_e1156, clk, rst, out_s1157, out_e1157, result1157);
PE P1158(out_s1094, out_e1157, clk, rst, out_s1158, out_e1158, result1158);
PE P1159(out_s1095, out_e1158, clk, rst, out_s1159, out_e1159, result1159);
PE P1160(out_s1096, out_e1159, clk, rst, out_s1160, out_e1160, result1160);
PE P1161(out_s1097, out_e1160, clk, rst, out_s1161, out_e1161, result1161);
PE P1162(out_s1098, out_e1161, clk, rst, out_s1162, out_e1162, result1162);
PE P1163(out_s1099, out_e1162, clk, rst, out_s1163, out_e1163, result1163);
PE P1164(out_s1100, out_e1163, clk, rst, out_s1164, out_e1164, result1164);
PE P1165(out_s1101, out_e1164, clk, rst, out_s1165, out_e1165, result1165);
PE P1166(out_s1102, out_e1165, clk, rst, out_s1166, out_e1166, result1166);
PE P1167(out_s1103, out_e1166, clk, rst, out_s1167, out_e1167, result1167);
PE P1168(out_s1104, out_e1167, clk, rst, out_s1168, out_e1168, result1168);
PE P1169(out_s1105, out_e1168, clk, rst, out_s1169, out_e1169, result1169);
PE P1170(out_s1106, out_e1169, clk, rst, out_s1170, out_e1170, result1170);
PE P1171(out_s1107, out_e1170, clk, rst, out_s1171, out_e1171, result1171);
PE P1172(out_s1108, out_e1171, clk, rst, out_s1172, out_e1172, result1172);
PE P1173(out_s1109, out_e1172, clk, rst, out_s1173, out_e1173, result1173);
PE P1174(out_s1110, out_e1173, clk, rst, out_s1174, out_e1174, result1174);
PE P1175(out_s1111, out_e1174, clk, rst, out_s1175, out_e1175, result1175);
PE P1176(out_s1112, out_e1175, clk, rst, out_s1176, out_e1176, result1176);
PE P1177(out_s1113, out_e1176, clk, rst, out_s1177, out_e1177, result1177);
PE P1178(out_s1114, out_e1177, clk, rst, out_s1178, out_e1178, result1178);
PE P1179(out_s1115, out_e1178, clk, rst, out_s1179, out_e1179, result1179);
PE P1180(out_s1116, out_e1179, clk, rst, out_s1180, out_e1180, result1180);
PE P1181(out_s1117, out_e1180, clk, rst, out_s1181, out_e1181, result1181);
PE P1182(out_s1118, out_e1181, clk, rst, out_s1182, out_e1182, result1182);
PE P1183(out_s1119, out_e1182, clk, rst, out_s1183, out_e1183, result1183);
PE P1184(out_s1120, out_e1183, clk, rst, out_s1184, out_e1184, result1184);
PE P1185(out_s1121, out_e1184, clk, rst, out_s1185, out_e1185, result1185);
PE P1186(out_s1122, out_e1185, clk, rst, out_s1186, out_e1186, result1186);
PE P1187(out_s1123, out_e1186, clk, rst, out_s1187, out_e1187, result1187);
PE P1188(out_s1124, out_e1187, clk, rst, out_s1188, out_e1188, result1188);
PE P1189(out_s1125, out_e1188, clk, rst, out_s1189, out_e1189, result1189);
PE P1190(out_s1126, out_e1189, clk, rst, out_s1190, out_e1190, result1190);
PE P1191(out_s1127, out_e1190, clk, rst, out_s1191, out_e1191, result1191);
PE P1192(out_s1128, out_e1191, clk, rst, out_s1192, out_e1192, result1192);
PE P1193(out_s1129, out_e1192, clk, rst, out_s1193, out_e1193, result1193);
PE P1194(out_s1130, out_e1193, clk, rst, out_s1194, out_e1194, result1194);
PE P1195(out_s1131, out_e1194, clk, rst, out_s1195, out_e1195, result1195);
PE P1196(out_s1132, out_e1195, clk, rst, out_s1196, out_e1196, result1196);
PE P1197(out_s1133, out_e1196, clk, rst, out_s1197, out_e1197, result1197);
PE P1198(out_s1134, out_e1197, clk, rst, out_s1198, out_e1198, result1198);
PE P1199(out_s1135, out_e1198, clk, rst, out_s1199, out_e1199, result1199);
PE P1200(out_s1136, out_e1199, clk, rst, out_s1200, out_e1200, result1200);
PE P1201(out_s1137, out_e1200, clk, rst, out_s1201, out_e1201, result1201);
PE P1202(out_s1138, out_e1201, clk, rst, out_s1202, out_e1202, result1202);
PE P1203(out_s1139, out_e1202, clk, rst, out_s1203, out_e1203, result1203);
PE P1204(out_s1140, out_e1203, clk, rst, out_s1204, out_e1204, result1204);
PE P1205(out_s1141, out_e1204, clk, rst, out_s1205, out_e1205, result1205);
PE P1206(out_s1142, out_e1205, clk, rst, out_s1206, out_e1206, result1206);
PE P1207(out_s1143, out_e1206, clk, rst, out_s1207, out_e1207, result1207);
PE P1208(out_s1144, out_e1207, clk, rst, out_s1208, out_e1208, result1208);
PE P1209(out_s1145, out_e1208, clk, rst, out_s1209, out_e1209, result1209);
PE P1210(out_s1146, out_e1209, clk, rst, out_s1210, out_e1210, result1210);
PE P1211(out_s1147, out_e1210, clk, rst, out_s1211, out_e1211, result1211);
PE P1212(out_s1148, out_e1211, clk, rst, out_s1212, out_e1212, result1212);
PE P1213(out_s1149, out_e1212, clk, rst, out_s1213, out_e1213, result1213);
PE P1214(out_s1150, out_e1213, clk, rst, out_s1214, out_e1214, result1214);
PE P1215(out_s1151, out_e1214, clk, rst, out_s1215, out_e1215, result1215);

PE P1217(out_s1153, out_e1216, clk, rst, out_s1217, out_e1217, result1217);
PE P1218(out_s1154, out_e1217, clk, rst, out_s1218, out_e1218, result1218);
PE P1219(out_s1155, out_e1218, clk, rst, out_s1219, out_e1219, result1219);
PE P1220(out_s1156, out_e1219, clk, rst, out_s1220, out_e1220, result1220);
PE P1221(out_s1157, out_e1220, clk, rst, out_s1221, out_e1221, result1221);
PE P1222(out_s1158, out_e1221, clk, rst, out_s1222, out_e1222, result1222);
PE P1223(out_s1159, out_e1222, clk, rst, out_s1223, out_e1223, result1223);
PE P1224(out_s1160, out_e1223, clk, rst, out_s1224, out_e1224, result1224);
PE P1225(out_s1161, out_e1224, clk, rst, out_s1225, out_e1225, result1225);
PE P1226(out_s1162, out_e1225, clk, rst, out_s1226, out_e1226, result1226);
PE P1227(out_s1163, out_e1226, clk, rst, out_s1227, out_e1227, result1227);
PE P1228(out_s1164, out_e1227, clk, rst, out_s1228, out_e1228, result1228);
PE P1229(out_s1165, out_e1228, clk, rst, out_s1229, out_e1229, result1229);
PE P1230(out_s1166, out_e1229, clk, rst, out_s1230, out_e1230, result1230);
PE P1231(out_s1167, out_e1230, clk, rst, out_s1231, out_e1231, result1231);
PE P1232(out_s1168, out_e1231, clk, rst, out_s1232, out_e1232, result1232);
PE P1233(out_s1169, out_e1232, clk, rst, out_s1233, out_e1233, result1233);
PE P1234(out_s1170, out_e1233, clk, rst, out_s1234, out_e1234, result1234);
PE P1235(out_s1171, out_e1234, clk, rst, out_s1235, out_e1235, result1235);
PE P1236(out_s1172, out_e1235, clk, rst, out_s1236, out_e1236, result1236);
PE P1237(out_s1173, out_e1236, clk, rst, out_s1237, out_e1237, result1237);
PE P1238(out_s1174, out_e1237, clk, rst, out_s1238, out_e1238, result1238);
PE P1239(out_s1175, out_e1238, clk, rst, out_s1239, out_e1239, result1239);
PE P1240(out_s1176, out_e1239, clk, rst, out_s1240, out_e1240, result1240);
PE P1241(out_s1177, out_e1240, clk, rst, out_s1241, out_e1241, result1241);
PE P1242(out_s1178, out_e1241, clk, rst, out_s1242, out_e1242, result1242);
PE P1243(out_s1179, out_e1242, clk, rst, out_s1243, out_e1243, result1243);
PE P1244(out_s1180, out_e1243, clk, rst, out_s1244, out_e1244, result1244);
PE P1245(out_s1181, out_e1244, clk, rst, out_s1245, out_e1245, result1245);
PE P1246(out_s1182, out_e1245, clk, rst, out_s1246, out_e1246, result1246);
PE P1247(out_s1183, out_e1246, clk, rst, out_s1247, out_e1247, result1247);
PE P1248(out_s1184, out_e1247, clk, rst, out_s1248, out_e1248, result1248);
PE P1249(out_s1185, out_e1248, clk, rst, out_s1249, out_e1249, result1249);
PE P1250(out_s1186, out_e1249, clk, rst, out_s1250, out_e1250, result1250);
PE P1251(out_s1187, out_e1250, clk, rst, out_s1251, out_e1251, result1251);
PE P1252(out_s1188, out_e1251, clk, rst, out_s1252, out_e1252, result1252);
PE P1253(out_s1189, out_e1252, clk, rst, out_s1253, out_e1253, result1253);
PE P1254(out_s1190, out_e1253, clk, rst, out_s1254, out_e1254, result1254);
PE P1255(out_s1191, out_e1254, clk, rst, out_s1255, out_e1255, result1255);
PE P1256(out_s1192, out_e1255, clk, rst, out_s1256, out_e1256, result1256);
PE P1257(out_s1193, out_e1256, clk, rst, out_s1257, out_e1257, result1257);
PE P1258(out_s1194, out_e1257, clk, rst, out_s1258, out_e1258, result1258);
PE P1259(out_s1195, out_e1258, clk, rst, out_s1259, out_e1259, result1259);
PE P1260(out_s1196, out_e1259, clk, rst, out_s1260, out_e1260, result1260);
PE P1261(out_s1197, out_e1260, clk, rst, out_s1261, out_e1261, result1261);
PE P1262(out_s1198, out_e1261, clk, rst, out_s1262, out_e1262, result1262);
PE P1263(out_s1199, out_e1262, clk, rst, out_s1263, out_e1263, result1263);
PE P1264(out_s1200, out_e1263, clk, rst, out_s1264, out_e1264, result1264);
PE P1265(out_s1201, out_e1264, clk, rst, out_s1265, out_e1265, result1265);
PE P1266(out_s1202, out_e1265, clk, rst, out_s1266, out_e1266, result1266);
PE P1267(out_s1203, out_e1266, clk, rst, out_s1267, out_e1267, result1267);
PE P1268(out_s1204, out_e1267, clk, rst, out_s1268, out_e1268, result1268);
PE P1269(out_s1205, out_e1268, clk, rst, out_s1269, out_e1269, result1269);
PE P1270(out_s1206, out_e1269, clk, rst, out_s1270, out_e1270, result1270);
PE P1271(out_s1207, out_e1270, clk, rst, out_s1271, out_e1271, result1271);
PE P1272(out_s1208, out_e1271, clk, rst, out_s1272, out_e1272, result1272);
PE P1273(out_s1209, out_e1272, clk, rst, out_s1273, out_e1273, result1273);
PE P1274(out_s1210, out_e1273, clk, rst, out_s1274, out_e1274, result1274);
PE P1275(out_s1211, out_e1274, clk, rst, out_s1275, out_e1275, result1275);
PE P1276(out_s1212, out_e1275, clk, rst, out_s1276, out_e1276, result1276);
PE P1277(out_s1213, out_e1276, clk, rst, out_s1277, out_e1277, result1277);
PE P1278(out_s1214, out_e1277, clk, rst, out_s1278, out_e1278, result1278);
PE P1279(out_s1215, out_e1278, clk, rst, out_s1279, out_e1279, result1279);

PE P1281(out_s1217, out_e1280, clk, rst, out_s1281, out_e1281, result1281);
PE P1282(out_s1218, out_e1281, clk, rst, out_s1282, out_e1282, result1282);
PE P1283(out_s1219, out_e1282, clk, rst, out_s1283, out_e1283, result1283);
PE P1284(out_s1220, out_e1283, clk, rst, out_s1284, out_e1284, result1284);
PE P1285(out_s1221, out_e1284, clk, rst, out_s1285, out_e1285, result1285);
PE P1286(out_s1222, out_e1285, clk, rst, out_s1286, out_e1286, result1286);
PE P1287(out_s1223, out_e1286, clk, rst, out_s1287, out_e1287, result1287);
PE P1288(out_s1224, out_e1287, clk, rst, out_s1288, out_e1288, result1288);
PE P1289(out_s1225, out_e1288, clk, rst, out_s1289, out_e1289, result1289);
PE P1290(out_s1226, out_e1289, clk, rst, out_s1290, out_e1290, result1290);
PE P1291(out_s1227, out_e1290, clk, rst, out_s1291, out_e1291, result1291);
PE P1292(out_s1228, out_e1291, clk, rst, out_s1292, out_e1292, result1292);
PE P1293(out_s1229, out_e1292, clk, rst, out_s1293, out_e1293, result1293);
PE P1294(out_s1230, out_e1293, clk, rst, out_s1294, out_e1294, result1294);
PE P1295(out_s1231, out_e1294, clk, rst, out_s1295, out_e1295, result1295);
PE P1296(out_s1232, out_e1295, clk, rst, out_s1296, out_e1296, result1296);
PE P1297(out_s1233, out_e1296, clk, rst, out_s1297, out_e1297, result1297);
PE P1298(out_s1234, out_e1297, clk, rst, out_s1298, out_e1298, result1298);
PE P1299(out_s1235, out_e1298, clk, rst, out_s1299, out_e1299, result1299);
PE P1300(out_s1236, out_e1299, clk, rst, out_s1300, out_e1300, result1300);
PE P1301(out_s1237, out_e1300, clk, rst, out_s1301, out_e1301, result1301);
PE P1302(out_s1238, out_e1301, clk, rst, out_s1302, out_e1302, result1302);
PE P1303(out_s1239, out_e1302, clk, rst, out_s1303, out_e1303, result1303);
PE P1304(out_s1240, out_e1303, clk, rst, out_s1304, out_e1304, result1304);
PE P1305(out_s1241, out_e1304, clk, rst, out_s1305, out_e1305, result1305);
PE P1306(out_s1242, out_e1305, clk, rst, out_s1306, out_e1306, result1306);
PE P1307(out_s1243, out_e1306, clk, rst, out_s1307, out_e1307, result1307);
PE P1308(out_s1244, out_e1307, clk, rst, out_s1308, out_e1308, result1308);
PE P1309(out_s1245, out_e1308, clk, rst, out_s1309, out_e1309, result1309);
PE P1310(out_s1246, out_e1309, clk, rst, out_s1310, out_e1310, result1310);
PE P1311(out_s1247, out_e1310, clk, rst, out_s1311, out_e1311, result1311);
PE P1312(out_s1248, out_e1311, clk, rst, out_s1312, out_e1312, result1312);
PE P1313(out_s1249, out_e1312, clk, rst, out_s1313, out_e1313, result1313);
PE P1314(out_s1250, out_e1313, clk, rst, out_s1314, out_e1314, result1314);
PE P1315(out_s1251, out_e1314, clk, rst, out_s1315, out_e1315, result1315);
PE P1316(out_s1252, out_e1315, clk, rst, out_s1316, out_e1316, result1316);
PE P1317(out_s1253, out_e1316, clk, rst, out_s1317, out_e1317, result1317);
PE P1318(out_s1254, out_e1317, clk, rst, out_s1318, out_e1318, result1318);
PE P1319(out_s1255, out_e1318, clk, rst, out_s1319, out_e1319, result1319);
PE P1320(out_s1256, out_e1319, clk, rst, out_s1320, out_e1320, result1320);
PE P1321(out_s1257, out_e1320, clk, rst, out_s1321, out_e1321, result1321);
PE P1322(out_s1258, out_e1321, clk, rst, out_s1322, out_e1322, result1322);
PE P1323(out_s1259, out_e1322, clk, rst, out_s1323, out_e1323, result1323);
PE P1324(out_s1260, out_e1323, clk, rst, out_s1324, out_e1324, result1324);
PE P1325(out_s1261, out_e1324, clk, rst, out_s1325, out_e1325, result1325);
PE P1326(out_s1262, out_e1325, clk, rst, out_s1326, out_e1326, result1326);
PE P1327(out_s1263, out_e1326, clk, rst, out_s1327, out_e1327, result1327);
PE P1328(out_s1264, out_e1327, clk, rst, out_s1328, out_e1328, result1328);
PE P1329(out_s1265, out_e1328, clk, rst, out_s1329, out_e1329, result1329);
PE P1330(out_s1266, out_e1329, clk, rst, out_s1330, out_e1330, result1330);
PE P1331(out_s1267, out_e1330, clk, rst, out_s1331, out_e1331, result1331);
PE P1332(out_s1268, out_e1331, clk, rst, out_s1332, out_e1332, result1332);
PE P1333(out_s1269, out_e1332, clk, rst, out_s1333, out_e1333, result1333);
PE P1334(out_s1270, out_e1333, clk, rst, out_s1334, out_e1334, result1334);
PE P1335(out_s1271, out_e1334, clk, rst, out_s1335, out_e1335, result1335);
PE P1336(out_s1272, out_e1335, clk, rst, out_s1336, out_e1336, result1336);
PE P1337(out_s1273, out_e1336, clk, rst, out_s1337, out_e1337, result1337);
PE P1338(out_s1274, out_e1337, clk, rst, out_s1338, out_e1338, result1338);
PE P1339(out_s1275, out_e1338, clk, rst, out_s1339, out_e1339, result1339);
PE P1340(out_s1276, out_e1339, clk, rst, out_s1340, out_e1340, result1340);
PE P1341(out_s1277, out_e1340, clk, rst, out_s1341, out_e1341, result1341);
PE P1342(out_s1278, out_e1341, clk, rst, out_s1342, out_e1342, result1342);
PE P1343(out_s1279, out_e1342, clk, rst, out_s1343, out_e1343, result1343);

PE P1345(out_s1281, out_e1344, clk, rst, out_s1345, out_e1345, result1345);
PE P1346(out_s1282, out_e1345, clk, rst, out_s1346, out_e1346, result1346);
PE P1347(out_s1283, out_e1346, clk, rst, out_s1347, out_e1347, result1347);
PE P1348(out_s1284, out_e1347, clk, rst, out_s1348, out_e1348, result1348);
PE P1349(out_s1285, out_e1348, clk, rst, out_s1349, out_e1349, result1349);
PE P1350(out_s1286, out_e1349, clk, rst, out_s1350, out_e1350, result1350);
PE P1351(out_s1287, out_e1350, clk, rst, out_s1351, out_e1351, result1351);
PE P1352(out_s1288, out_e1351, clk, rst, out_s1352, out_e1352, result1352);
PE P1353(out_s1289, out_e1352, clk, rst, out_s1353, out_e1353, result1353);
PE P1354(out_s1290, out_e1353, clk, rst, out_s1354, out_e1354, result1354);
PE P1355(out_s1291, out_e1354, clk, rst, out_s1355, out_e1355, result1355);
PE P1356(out_s1292, out_e1355, clk, rst, out_s1356, out_e1356, result1356);
PE P1357(out_s1293, out_e1356, clk, rst, out_s1357, out_e1357, result1357);
PE P1358(out_s1294, out_e1357, clk, rst, out_s1358, out_e1358, result1358);
PE P1359(out_s1295, out_e1358, clk, rst, out_s1359, out_e1359, result1359);
PE P1360(out_s1296, out_e1359, clk, rst, out_s1360, out_e1360, result1360);
PE P1361(out_s1297, out_e1360, clk, rst, out_s1361, out_e1361, result1361);
PE P1362(out_s1298, out_e1361, clk, rst, out_s1362, out_e1362, result1362);
PE P1363(out_s1299, out_e1362, clk, rst, out_s1363, out_e1363, result1363);
PE P1364(out_s1300, out_e1363, clk, rst, out_s1364, out_e1364, result1364);
PE P1365(out_s1301, out_e1364, clk, rst, out_s1365, out_e1365, result1365);
PE P1366(out_s1302, out_e1365, clk, rst, out_s1366, out_e1366, result1366);
PE P1367(out_s1303, out_e1366, clk, rst, out_s1367, out_e1367, result1367);
PE P1368(out_s1304, out_e1367, clk, rst, out_s1368, out_e1368, result1368);
PE P1369(out_s1305, out_e1368, clk, rst, out_s1369, out_e1369, result1369);
PE P1370(out_s1306, out_e1369, clk, rst, out_s1370, out_e1370, result1370);
PE P1371(out_s1307, out_e1370, clk, rst, out_s1371, out_e1371, result1371);
PE P1372(out_s1308, out_e1371, clk, rst, out_s1372, out_e1372, result1372);
PE P1373(out_s1309, out_e1372, clk, rst, out_s1373, out_e1373, result1373);
PE P1374(out_s1310, out_e1373, clk, rst, out_s1374, out_e1374, result1374);
PE P1375(out_s1311, out_e1374, clk, rst, out_s1375, out_e1375, result1375);
PE P1376(out_s1312, out_e1375, clk, rst, out_s1376, out_e1376, result1376);
PE P1377(out_s1313, out_e1376, clk, rst, out_s1377, out_e1377, result1377);
PE P1378(out_s1314, out_e1377, clk, rst, out_s1378, out_e1378, result1378);
PE P1379(out_s1315, out_e1378, clk, rst, out_s1379, out_e1379, result1379);
PE P1380(out_s1316, out_e1379, clk, rst, out_s1380, out_e1380, result1380);
PE P1381(out_s1317, out_e1380, clk, rst, out_s1381, out_e1381, result1381);
PE P1382(out_s1318, out_e1381, clk, rst, out_s1382, out_e1382, result1382);
PE P1383(out_s1319, out_e1382, clk, rst, out_s1383, out_e1383, result1383);
PE P1384(out_s1320, out_e1383, clk, rst, out_s1384, out_e1384, result1384);
PE P1385(out_s1321, out_e1384, clk, rst, out_s1385, out_e1385, result1385);
PE P1386(out_s1322, out_e1385, clk, rst, out_s1386, out_e1386, result1386);
PE P1387(out_s1323, out_e1386, clk, rst, out_s1387, out_e1387, result1387);
PE P1388(out_s1324, out_e1387, clk, rst, out_s1388, out_e1388, result1388);
PE P1389(out_s1325, out_e1388, clk, rst, out_s1389, out_e1389, result1389);
PE P1390(out_s1326, out_e1389, clk, rst, out_s1390, out_e1390, result1390);
PE P1391(out_s1327, out_e1390, clk, rst, out_s1391, out_e1391, result1391);
PE P1392(out_s1328, out_e1391, clk, rst, out_s1392, out_e1392, result1392);
PE P1393(out_s1329, out_e1392, clk, rst, out_s1393, out_e1393, result1393);
PE P1394(out_s1330, out_e1393, clk, rst, out_s1394, out_e1394, result1394);
PE P1395(out_s1331, out_e1394, clk, rst, out_s1395, out_e1395, result1395);
PE P1396(out_s1332, out_e1395, clk, rst, out_s1396, out_e1396, result1396);
PE P1397(out_s1333, out_e1396, clk, rst, out_s1397, out_e1397, result1397);
PE P1398(out_s1334, out_e1397, clk, rst, out_s1398, out_e1398, result1398);
PE P1399(out_s1335, out_e1398, clk, rst, out_s1399, out_e1399, result1399);
PE P1400(out_s1336, out_e1399, clk, rst, out_s1400, out_e1400, result1400);
PE P1401(out_s1337, out_e1400, clk, rst, out_s1401, out_e1401, result1401);
PE P1402(out_s1338, out_e1401, clk, rst, out_s1402, out_e1402, result1402);
PE P1403(out_s1339, out_e1402, clk, rst, out_s1403, out_e1403, result1403);
PE P1404(out_s1340, out_e1403, clk, rst, out_s1404, out_e1404, result1404);
PE P1405(out_s1341, out_e1404, clk, rst, out_s1405, out_e1405, result1405);
PE P1406(out_s1342, out_e1405, clk, rst, out_s1406, out_e1406, result1406);
PE P1407(out_s1343, out_e1406, clk, rst, out_s1407, out_e1407, result1407);

PE P1409(out_s1345, out_e1408, clk, rst, out_s1409, out_e1409, result1409);
PE P1410(out_s1346, out_e1409, clk, rst, out_s1410, out_e1410, result1410);
PE P1411(out_s1347, out_e1410, clk, rst, out_s1411, out_e1411, result1411);
PE P1412(out_s1348, out_e1411, clk, rst, out_s1412, out_e1412, result1412);
PE P1413(out_s1349, out_e1412, clk, rst, out_s1413, out_e1413, result1413);
PE P1414(out_s1350, out_e1413, clk, rst, out_s1414, out_e1414, result1414);
PE P1415(out_s1351, out_e1414, clk, rst, out_s1415, out_e1415, result1415);
PE P1416(out_s1352, out_e1415, clk, rst, out_s1416, out_e1416, result1416);
PE P1417(out_s1353, out_e1416, clk, rst, out_s1417, out_e1417, result1417);
PE P1418(out_s1354, out_e1417, clk, rst, out_s1418, out_e1418, result1418);
PE P1419(out_s1355, out_e1418, clk, rst, out_s1419, out_e1419, result1419);
PE P1420(out_s1356, out_e1419, clk, rst, out_s1420, out_e1420, result1420);
PE P1421(out_s1357, out_e1420, clk, rst, out_s1421, out_e1421, result1421);
PE P1422(out_s1358, out_e1421, clk, rst, out_s1422, out_e1422, result1422);
PE P1423(out_s1359, out_e1422, clk, rst, out_s1423, out_e1423, result1423);
PE P1424(out_s1360, out_e1423, clk, rst, out_s1424, out_e1424, result1424);
PE P1425(out_s1361, out_e1424, clk, rst, out_s1425, out_e1425, result1425);
PE P1426(out_s1362, out_e1425, clk, rst, out_s1426, out_e1426, result1426);
PE P1427(out_s1363, out_e1426, clk, rst, out_s1427, out_e1427, result1427);
PE P1428(out_s1364, out_e1427, clk, rst, out_s1428, out_e1428, result1428);
PE P1429(out_s1365, out_e1428, clk, rst, out_s1429, out_e1429, result1429);
PE P1430(out_s1366, out_e1429, clk, rst, out_s1430, out_e1430, result1430);
PE P1431(out_s1367, out_e1430, clk, rst, out_s1431, out_e1431, result1431);
PE P1432(out_s1368, out_e1431, clk, rst, out_s1432, out_e1432, result1432);
PE P1433(out_s1369, out_e1432, clk, rst, out_s1433, out_e1433, result1433);
PE P1434(out_s1370, out_e1433, clk, rst, out_s1434, out_e1434, result1434);
PE P1435(out_s1371, out_e1434, clk, rst, out_s1435, out_e1435, result1435);
PE P1436(out_s1372, out_e1435, clk, rst, out_s1436, out_e1436, result1436);
PE P1437(out_s1373, out_e1436, clk, rst, out_s1437, out_e1437, result1437);
PE P1438(out_s1374, out_e1437, clk, rst, out_s1438, out_e1438, result1438);
PE P1439(out_s1375, out_e1438, clk, rst, out_s1439, out_e1439, result1439);
PE P1440(out_s1376, out_e1439, clk, rst, out_s1440, out_e1440, result1440);
PE P1441(out_s1377, out_e1440, clk, rst, out_s1441, out_e1441, result1441);
PE P1442(out_s1378, out_e1441, clk, rst, out_s1442, out_e1442, result1442);
PE P1443(out_s1379, out_e1442, clk, rst, out_s1443, out_e1443, result1443);
PE P1444(out_s1380, out_e1443, clk, rst, out_s1444, out_e1444, result1444);
PE P1445(out_s1381, out_e1444, clk, rst, out_s1445, out_e1445, result1445);
PE P1446(out_s1382, out_e1445, clk, rst, out_s1446, out_e1446, result1446);
PE P1447(out_s1383, out_e1446, clk, rst, out_s1447, out_e1447, result1447);
PE P1448(out_s1384, out_e1447, clk, rst, out_s1448, out_e1448, result1448);
PE P1449(out_s1385, out_e1448, clk, rst, out_s1449, out_e1449, result1449);
PE P1450(out_s1386, out_e1449, clk, rst, out_s1450, out_e1450, result1450);
PE P1451(out_s1387, out_e1450, clk, rst, out_s1451, out_e1451, result1451);
PE P1452(out_s1388, out_e1451, clk, rst, out_s1452, out_e1452, result1452);
PE P1453(out_s1389, out_e1452, clk, rst, out_s1453, out_e1453, result1453);
PE P1454(out_s1390, out_e1453, clk, rst, out_s1454, out_e1454, result1454);
PE P1455(out_s1391, out_e1454, clk, rst, out_s1455, out_e1455, result1455);
PE P1456(out_s1392, out_e1455, clk, rst, out_s1456, out_e1456, result1456);
PE P1457(out_s1393, out_e1456, clk, rst, out_s1457, out_e1457, result1457);
PE P1458(out_s1394, out_e1457, clk, rst, out_s1458, out_e1458, result1458);
PE P1459(out_s1395, out_e1458, clk, rst, out_s1459, out_e1459, result1459);
PE P1460(out_s1396, out_e1459, clk, rst, out_s1460, out_e1460, result1460);
PE P1461(out_s1397, out_e1460, clk, rst, out_s1461, out_e1461, result1461);
PE P1462(out_s1398, out_e1461, clk, rst, out_s1462, out_e1462, result1462);
PE P1463(out_s1399, out_e1462, clk, rst, out_s1463, out_e1463, result1463);
PE P1464(out_s1400, out_e1463, clk, rst, out_s1464, out_e1464, result1464);
PE P1465(out_s1401, out_e1464, clk, rst, out_s1465, out_e1465, result1465);
PE P1466(out_s1402, out_e1465, clk, rst, out_s1466, out_e1466, result1466);
PE P1467(out_s1403, out_e1466, clk, rst, out_s1467, out_e1467, result1467);
PE P1468(out_s1404, out_e1467, clk, rst, out_s1468, out_e1468, result1468);
PE P1469(out_s1405, out_e1468, clk, rst, out_s1469, out_e1469, result1469);
PE P1470(out_s1406, out_e1469, clk, rst, out_s1470, out_e1470, result1470);
PE P1471(out_s1407, out_e1470, clk, rst, out_s1471, out_e1471, result1471);

PE P1473(out_s1409, out_e1472, clk, rst, out_s1473, out_e1473, result1473);
PE P1474(out_s1410, out_e1473, clk, rst, out_s1474, out_e1474, result1474);
PE P1475(out_s1411, out_e1474, clk, rst, out_s1475, out_e1475, result1475);
PE P1476(out_s1412, out_e1475, clk, rst, out_s1476, out_e1476, result1476);
PE P1477(out_s1413, out_e1476, clk, rst, out_s1477, out_e1477, result1477);
PE P1478(out_s1414, out_e1477, clk, rst, out_s1478, out_e1478, result1478);
PE P1479(out_s1415, out_e1478, clk, rst, out_s1479, out_e1479, result1479);
PE P1480(out_s1416, out_e1479, clk, rst, out_s1480, out_e1480, result1480);
PE P1481(out_s1417, out_e1480, clk, rst, out_s1481, out_e1481, result1481);
PE P1482(out_s1418, out_e1481, clk, rst, out_s1482, out_e1482, result1482);
PE P1483(out_s1419, out_e1482, clk, rst, out_s1483, out_e1483, result1483);
PE P1484(out_s1420, out_e1483, clk, rst, out_s1484, out_e1484, result1484);
PE P1485(out_s1421, out_e1484, clk, rst, out_s1485, out_e1485, result1485);
PE P1486(out_s1422, out_e1485, clk, rst, out_s1486, out_e1486, result1486);
PE P1487(out_s1423, out_e1486, clk, rst, out_s1487, out_e1487, result1487);
PE P1488(out_s1424, out_e1487, clk, rst, out_s1488, out_e1488, result1488);
PE P1489(out_s1425, out_e1488, clk, rst, out_s1489, out_e1489, result1489);
PE P1490(out_s1426, out_e1489, clk, rst, out_s1490, out_e1490, result1490);
PE P1491(out_s1427, out_e1490, clk, rst, out_s1491, out_e1491, result1491);
PE P1492(out_s1428, out_e1491, clk, rst, out_s1492, out_e1492, result1492);
PE P1493(out_s1429, out_e1492, clk, rst, out_s1493, out_e1493, result1493);
PE P1494(out_s1430, out_e1493, clk, rst, out_s1494, out_e1494, result1494);
PE P1495(out_s1431, out_e1494, clk, rst, out_s1495, out_e1495, result1495);
PE P1496(out_s1432, out_e1495, clk, rst, out_s1496, out_e1496, result1496);
PE P1497(out_s1433, out_e1496, clk, rst, out_s1497, out_e1497, result1497);
PE P1498(out_s1434, out_e1497, clk, rst, out_s1498, out_e1498, result1498);
PE P1499(out_s1435, out_e1498, clk, rst, out_s1499, out_e1499, result1499);
PE P1500(out_s1436, out_e1499, clk, rst, out_s1500, out_e1500, result1500);
PE P1501(out_s1437, out_e1500, clk, rst, out_s1501, out_e1501, result1501);
PE P1502(out_s1438, out_e1501, clk, rst, out_s1502, out_e1502, result1502);
PE P1503(out_s1439, out_e1502, clk, rst, out_s1503, out_e1503, result1503);
PE P1504(out_s1440, out_e1503, clk, rst, out_s1504, out_e1504, result1504);
PE P1505(out_s1441, out_e1504, clk, rst, out_s1505, out_e1505, result1505);
PE P1506(out_s1442, out_e1505, clk, rst, out_s1506, out_e1506, result1506);
PE P1507(out_s1443, out_e1506, clk, rst, out_s1507, out_e1507, result1507);
PE P1508(out_s1444, out_e1507, clk, rst, out_s1508, out_e1508, result1508);
PE P1509(out_s1445, out_e1508, clk, rst, out_s1509, out_e1509, result1509);
PE P1510(out_s1446, out_e1509, clk, rst, out_s1510, out_e1510, result1510);
PE P1511(out_s1447, out_e1510, clk, rst, out_s1511, out_e1511, result1511);
PE P1512(out_s1448, out_e1511, clk, rst, out_s1512, out_e1512, result1512);
PE P1513(out_s1449, out_e1512, clk, rst, out_s1513, out_e1513, result1513);
PE P1514(out_s1450, out_e1513, clk, rst, out_s1514, out_e1514, result1514);
PE P1515(out_s1451, out_e1514, clk, rst, out_s1515, out_e1515, result1515);
PE P1516(out_s1452, out_e1515, clk, rst, out_s1516, out_e1516, result1516);
PE P1517(out_s1453, out_e1516, clk, rst, out_s1517, out_e1517, result1517);
PE P1518(out_s1454, out_e1517, clk, rst, out_s1518, out_e1518, result1518);
PE P1519(out_s1455, out_e1518, clk, rst, out_s1519, out_e1519, result1519);
PE P1520(out_s1456, out_e1519, clk, rst, out_s1520, out_e1520, result1520);
PE P1521(out_s1457, out_e1520, clk, rst, out_s1521, out_e1521, result1521);
PE P1522(out_s1458, out_e1521, clk, rst, out_s1522, out_e1522, result1522);
PE P1523(out_s1459, out_e1522, clk, rst, out_s1523, out_e1523, result1523);
PE P1524(out_s1460, out_e1523, clk, rst, out_s1524, out_e1524, result1524);
PE P1525(out_s1461, out_e1524, clk, rst, out_s1525, out_e1525, result1525);
PE P1526(out_s1462, out_e1525, clk, rst, out_s1526, out_e1526, result1526);
PE P1527(out_s1463, out_e1526, clk, rst, out_s1527, out_e1527, result1527);
PE P1528(out_s1464, out_e1527, clk, rst, out_s1528, out_e1528, result1528);
PE P1529(out_s1465, out_e1528, clk, rst, out_s1529, out_e1529, result1529);
PE P1530(out_s1466, out_e1529, clk, rst, out_s1530, out_e1530, result1530);
PE P1531(out_s1467, out_e1530, clk, rst, out_s1531, out_e1531, result1531);
PE P1532(out_s1468, out_e1531, clk, rst, out_s1532, out_e1532, result1532);
PE P1533(out_s1469, out_e1532, clk, rst, out_s1533, out_e1533, result1533);
PE P1534(out_s1470, out_e1533, clk, rst, out_s1534, out_e1534, result1534);
PE P1535(out_s1471, out_e1534, clk, rst, out_s1535, out_e1535, result1535);

PE P1537(out_s1473, out_e1536, clk, rst, out_s1537, out_e1537, result1537);
PE P1538(out_s1474, out_e1537, clk, rst, out_s1538, out_e1538, result1538);
PE P1539(out_s1475, out_e1538, clk, rst, out_s1539, out_e1539, result1539);
PE P1540(out_s1476, out_e1539, clk, rst, out_s1540, out_e1540, result1540);
PE P1541(out_s1477, out_e1540, clk, rst, out_s1541, out_e1541, result1541);
PE P1542(out_s1478, out_e1541, clk, rst, out_s1542, out_e1542, result1542);
PE P1543(out_s1479, out_e1542, clk, rst, out_s1543, out_e1543, result1543);
PE P1544(out_s1480, out_e1543, clk, rst, out_s1544, out_e1544, result1544);
PE P1545(out_s1481, out_e1544, clk, rst, out_s1545, out_e1545, result1545);
PE P1546(out_s1482, out_e1545, clk, rst, out_s1546, out_e1546, result1546);
PE P1547(out_s1483, out_e1546, clk, rst, out_s1547, out_e1547, result1547);
PE P1548(out_s1484, out_e1547, clk, rst, out_s1548, out_e1548, result1548);
PE P1549(out_s1485, out_e1548, clk, rst, out_s1549, out_e1549, result1549);
PE P1550(out_s1486, out_e1549, clk, rst, out_s1550, out_e1550, result1550);
PE P1551(out_s1487, out_e1550, clk, rst, out_s1551, out_e1551, result1551);
PE P1552(out_s1488, out_e1551, clk, rst, out_s1552, out_e1552, result1552);
PE P1553(out_s1489, out_e1552, clk, rst, out_s1553, out_e1553, result1553);
PE P1554(out_s1490, out_e1553, clk, rst, out_s1554, out_e1554, result1554);
PE P1555(out_s1491, out_e1554, clk, rst, out_s1555, out_e1555, result1555);
PE P1556(out_s1492, out_e1555, clk, rst, out_s1556, out_e1556, result1556);
PE P1557(out_s1493, out_e1556, clk, rst, out_s1557, out_e1557, result1557);
PE P1558(out_s1494, out_e1557, clk, rst, out_s1558, out_e1558, result1558);
PE P1559(out_s1495, out_e1558, clk, rst, out_s1559, out_e1559, result1559);
PE P1560(out_s1496, out_e1559, clk, rst, out_s1560, out_e1560, result1560);
PE P1561(out_s1497, out_e1560, clk, rst, out_s1561, out_e1561, result1561);
PE P1562(out_s1498, out_e1561, clk, rst, out_s1562, out_e1562, result1562);
PE P1563(out_s1499, out_e1562, clk, rst, out_s1563, out_e1563, result1563);
PE P1564(out_s1500, out_e1563, clk, rst, out_s1564, out_e1564, result1564);
PE P1565(out_s1501, out_e1564, clk, rst, out_s1565, out_e1565, result1565);
PE P1566(out_s1502, out_e1565, clk, rst, out_s1566, out_e1566, result1566);
PE P1567(out_s1503, out_e1566, clk, rst, out_s1567, out_e1567, result1567);
PE P1568(out_s1504, out_e1567, clk, rst, out_s1568, out_e1568, result1568);
PE P1569(out_s1505, out_e1568, clk, rst, out_s1569, out_e1569, result1569);
PE P1570(out_s1506, out_e1569, clk, rst, out_s1570, out_e1570, result1570);
PE P1571(out_s1507, out_e1570, clk, rst, out_s1571, out_e1571, result1571);
PE P1572(out_s1508, out_e1571, clk, rst, out_s1572, out_e1572, result1572);
PE P1573(out_s1509, out_e1572, clk, rst, out_s1573, out_e1573, result1573);
PE P1574(out_s1510, out_e1573, clk, rst, out_s1574, out_e1574, result1574);
PE P1575(out_s1511, out_e1574, clk, rst, out_s1575, out_e1575, result1575);
PE P1576(out_s1512, out_e1575, clk, rst, out_s1576, out_e1576, result1576);
PE P1577(out_s1513, out_e1576, clk, rst, out_s1577, out_e1577, result1577);
PE P1578(out_s1514, out_e1577, clk, rst, out_s1578, out_e1578, result1578);
PE P1579(out_s1515, out_e1578, clk, rst, out_s1579, out_e1579, result1579);
PE P1580(out_s1516, out_e1579, clk, rst, out_s1580, out_e1580, result1580);
PE P1581(out_s1517, out_e1580, clk, rst, out_s1581, out_e1581, result1581);
PE P1582(out_s1518, out_e1581, clk, rst, out_s1582, out_e1582, result1582);
PE P1583(out_s1519, out_e1582, clk, rst, out_s1583, out_e1583, result1583);
PE P1584(out_s1520, out_e1583, clk, rst, out_s1584, out_e1584, result1584);
PE P1585(out_s1521, out_e1584, clk, rst, out_s1585, out_e1585, result1585);
PE P1586(out_s1522, out_e1585, clk, rst, out_s1586, out_e1586, result1586);
PE P1587(out_s1523, out_e1586, clk, rst, out_s1587, out_e1587, result1587);
PE P1588(out_s1524, out_e1587, clk, rst, out_s1588, out_e1588, result1588);
PE P1589(out_s1525, out_e1588, clk, rst, out_s1589, out_e1589, result1589);
PE P1590(out_s1526, out_e1589, clk, rst, out_s1590, out_e1590, result1590);
PE P1591(out_s1527, out_e1590, clk, rst, out_s1591, out_e1591, result1591);
PE P1592(out_s1528, out_e1591, clk, rst, out_s1592, out_e1592, result1592);
PE P1593(out_s1529, out_e1592, clk, rst, out_s1593, out_e1593, result1593);
PE P1594(out_s1530, out_e1593, clk, rst, out_s1594, out_e1594, result1594);
PE P1595(out_s1531, out_e1594, clk, rst, out_s1595, out_e1595, result1595);
PE P1596(out_s1532, out_e1595, clk, rst, out_s1596, out_e1596, result1596);
PE P1597(out_s1533, out_e1596, clk, rst, out_s1597, out_e1597, result1597);
PE P1598(out_s1534, out_e1597, clk, rst, out_s1598, out_e1598, result1598);
PE P1599(out_s1535, out_e1598, clk, rst, out_s1599, out_e1599, result1599);

PE P1601(out_s1537, out_e1600, clk, rst, out_s1601, out_e1601, result1601);
PE P1602(out_s1538, out_e1601, clk, rst, out_s1602, out_e1602, result1602);
PE P1603(out_s1539, out_e1602, clk, rst, out_s1603, out_e1603, result1603);
PE P1604(out_s1540, out_e1603, clk, rst, out_s1604, out_e1604, result1604);
PE P1605(out_s1541, out_e1604, clk, rst, out_s1605, out_e1605, result1605);
PE P1606(out_s1542, out_e1605, clk, rst, out_s1606, out_e1606, result1606);
PE P1607(out_s1543, out_e1606, clk, rst, out_s1607, out_e1607, result1607);
PE P1608(out_s1544, out_e1607, clk, rst, out_s1608, out_e1608, result1608);
PE P1609(out_s1545, out_e1608, clk, rst, out_s1609, out_e1609, result1609);
PE P1610(out_s1546, out_e1609, clk, rst, out_s1610, out_e1610, result1610);
PE P1611(out_s1547, out_e1610, clk, rst, out_s1611, out_e1611, result1611);
PE P1612(out_s1548, out_e1611, clk, rst, out_s1612, out_e1612, result1612);
PE P1613(out_s1549, out_e1612, clk, rst, out_s1613, out_e1613, result1613);
PE P1614(out_s1550, out_e1613, clk, rst, out_s1614, out_e1614, result1614);
PE P1615(out_s1551, out_e1614, clk, rst, out_s1615, out_e1615, result1615);
PE P1616(out_s1552, out_e1615, clk, rst, out_s1616, out_e1616, result1616);
PE P1617(out_s1553, out_e1616, clk, rst, out_s1617, out_e1617, result1617);
PE P1618(out_s1554, out_e1617, clk, rst, out_s1618, out_e1618, result1618);
PE P1619(out_s1555, out_e1618, clk, rst, out_s1619, out_e1619, result1619);
PE P1620(out_s1556, out_e1619, clk, rst, out_s1620, out_e1620, result1620);
PE P1621(out_s1557, out_e1620, clk, rst, out_s1621, out_e1621, result1621);
PE P1622(out_s1558, out_e1621, clk, rst, out_s1622, out_e1622, result1622);
PE P1623(out_s1559, out_e1622, clk, rst, out_s1623, out_e1623, result1623);
PE P1624(out_s1560, out_e1623, clk, rst, out_s1624, out_e1624, result1624);
PE P1625(out_s1561, out_e1624, clk, rst, out_s1625, out_e1625, result1625);
PE P1626(out_s1562, out_e1625, clk, rst, out_s1626, out_e1626, result1626);
PE P1627(out_s1563, out_e1626, clk, rst, out_s1627, out_e1627, result1627);
PE P1628(out_s1564, out_e1627, clk, rst, out_s1628, out_e1628, result1628);
PE P1629(out_s1565, out_e1628, clk, rst, out_s1629, out_e1629, result1629);
PE P1630(out_s1566, out_e1629, clk, rst, out_s1630, out_e1630, result1630);
PE P1631(out_s1567, out_e1630, clk, rst, out_s1631, out_e1631, result1631);
PE P1632(out_s1568, out_e1631, clk, rst, out_s1632, out_e1632, result1632);
PE P1633(out_s1569, out_e1632, clk, rst, out_s1633, out_e1633, result1633);
PE P1634(out_s1570, out_e1633, clk, rst, out_s1634, out_e1634, result1634);
PE P1635(out_s1571, out_e1634, clk, rst, out_s1635, out_e1635, result1635);
PE P1636(out_s1572, out_e1635, clk, rst, out_s1636, out_e1636, result1636);
PE P1637(out_s1573, out_e1636, clk, rst, out_s1637, out_e1637, result1637);
PE P1638(out_s1574, out_e1637, clk, rst, out_s1638, out_e1638, result1638);
PE P1639(out_s1575, out_e1638, clk, rst, out_s1639, out_e1639, result1639);
PE P1640(out_s1576, out_e1639, clk, rst, out_s1640, out_e1640, result1640);
PE P1641(out_s1577, out_e1640, clk, rst, out_s1641, out_e1641, result1641);
PE P1642(out_s1578, out_e1641, clk, rst, out_s1642, out_e1642, result1642);
PE P1643(out_s1579, out_e1642, clk, rst, out_s1643, out_e1643, result1643);
PE P1644(out_s1580, out_e1643, clk, rst, out_s1644, out_e1644, result1644);
PE P1645(out_s1581, out_e1644, clk, rst, out_s1645, out_e1645, result1645);
PE P1646(out_s1582, out_e1645, clk, rst, out_s1646, out_e1646, result1646);
PE P1647(out_s1583, out_e1646, clk, rst, out_s1647, out_e1647, result1647);
PE P1648(out_s1584, out_e1647, clk, rst, out_s1648, out_e1648, result1648);
PE P1649(out_s1585, out_e1648, clk, rst, out_s1649, out_e1649, result1649);
PE P1650(out_s1586, out_e1649, clk, rst, out_s1650, out_e1650, result1650);
PE P1651(out_s1587, out_e1650, clk, rst, out_s1651, out_e1651, result1651);
PE P1652(out_s1588, out_e1651, clk, rst, out_s1652, out_e1652, result1652);
PE P1653(out_s1589, out_e1652, clk, rst, out_s1653, out_e1653, result1653);
PE P1654(out_s1590, out_e1653, clk, rst, out_s1654, out_e1654, result1654);
PE P1655(out_s1591, out_e1654, clk, rst, out_s1655, out_e1655, result1655);
PE P1656(out_s1592, out_e1655, clk, rst, out_s1656, out_e1656, result1656);
PE P1657(out_s1593, out_e1656, clk, rst, out_s1657, out_e1657, result1657);
PE P1658(out_s1594, out_e1657, clk, rst, out_s1658, out_e1658, result1658);
PE P1659(out_s1595, out_e1658, clk, rst, out_s1659, out_e1659, result1659);
PE P1660(out_s1596, out_e1659, clk, rst, out_s1660, out_e1660, result1660);
PE P1661(out_s1597, out_e1660, clk, rst, out_s1661, out_e1661, result1661);
PE P1662(out_s1598, out_e1661, clk, rst, out_s1662, out_e1662, result1662);
PE P1663(out_s1599, out_e1662, clk, rst, out_s1663, out_e1663, result1663);

PE P1665(out_s1601, out_e1664, clk, rst, out_s1665, out_e1665, result1665);
PE P1666(out_s1602, out_e1665, clk, rst, out_s1666, out_e1666, result1666);
PE P1667(out_s1603, out_e1666, clk, rst, out_s1667, out_e1667, result1667);
PE P1668(out_s1604, out_e1667, clk, rst, out_s1668, out_e1668, result1668);
PE P1669(out_s1605, out_e1668, clk, rst, out_s1669, out_e1669, result1669);
PE P1670(out_s1606, out_e1669, clk, rst, out_s1670, out_e1670, result1670);
PE P1671(out_s1607, out_e1670, clk, rst, out_s1671, out_e1671, result1671);
PE P1672(out_s1608, out_e1671, clk, rst, out_s1672, out_e1672, result1672);
PE P1673(out_s1609, out_e1672, clk, rst, out_s1673, out_e1673, result1673);
PE P1674(out_s1610, out_e1673, clk, rst, out_s1674, out_e1674, result1674);
PE P1675(out_s1611, out_e1674, clk, rst, out_s1675, out_e1675, result1675);
PE P1676(out_s1612, out_e1675, clk, rst, out_s1676, out_e1676, result1676);
PE P1677(out_s1613, out_e1676, clk, rst, out_s1677, out_e1677, result1677);
PE P1678(out_s1614, out_e1677, clk, rst, out_s1678, out_e1678, result1678);
PE P1679(out_s1615, out_e1678, clk, rst, out_s1679, out_e1679, result1679);
PE P1680(out_s1616, out_e1679, clk, rst, out_s1680, out_e1680, result1680);
PE P1681(out_s1617, out_e1680, clk, rst, out_s1681, out_e1681, result1681);
PE P1682(out_s1618, out_e1681, clk, rst, out_s1682, out_e1682, result1682);
PE P1683(out_s1619, out_e1682, clk, rst, out_s1683, out_e1683, result1683);
PE P1684(out_s1620, out_e1683, clk, rst, out_s1684, out_e1684, result1684);
PE P1685(out_s1621, out_e1684, clk, rst, out_s1685, out_e1685, result1685);
PE P1686(out_s1622, out_e1685, clk, rst, out_s1686, out_e1686, result1686);
PE P1687(out_s1623, out_e1686, clk, rst, out_s1687, out_e1687, result1687);
PE P1688(out_s1624, out_e1687, clk, rst, out_s1688, out_e1688, result1688);
PE P1689(out_s1625, out_e1688, clk, rst, out_s1689, out_e1689, result1689);
PE P1690(out_s1626, out_e1689, clk, rst, out_s1690, out_e1690, result1690);
PE P1691(out_s1627, out_e1690, clk, rst, out_s1691, out_e1691, result1691);
PE P1692(out_s1628, out_e1691, clk, rst, out_s1692, out_e1692, result1692);
PE P1693(out_s1629, out_e1692, clk, rst, out_s1693, out_e1693, result1693);
PE P1694(out_s1630, out_e1693, clk, rst, out_s1694, out_e1694, result1694);
PE P1695(out_s1631, out_e1694, clk, rst, out_s1695, out_e1695, result1695);
PE P1696(out_s1632, out_e1695, clk, rst, out_s1696, out_e1696, result1696);
PE P1697(out_s1633, out_e1696, clk, rst, out_s1697, out_e1697, result1697);
PE P1698(out_s1634, out_e1697, clk, rst, out_s1698, out_e1698, result1698);
PE P1699(out_s1635, out_e1698, clk, rst, out_s1699, out_e1699, result1699);
PE P1700(out_s1636, out_e1699, clk, rst, out_s1700, out_e1700, result1700);
PE P1701(out_s1637, out_e1700, clk, rst, out_s1701, out_e1701, result1701);
PE P1702(out_s1638, out_e1701, clk, rst, out_s1702, out_e1702, result1702);
PE P1703(out_s1639, out_e1702, clk, rst, out_s1703, out_e1703, result1703);
PE P1704(out_s1640, out_e1703, clk, rst, out_s1704, out_e1704, result1704);
PE P1705(out_s1641, out_e1704, clk, rst, out_s1705, out_e1705, result1705);
PE P1706(out_s1642, out_e1705, clk, rst, out_s1706, out_e1706, result1706);
PE P1707(out_s1643, out_e1706, clk, rst, out_s1707, out_e1707, result1707);
PE P1708(out_s1644, out_e1707, clk, rst, out_s1708, out_e1708, result1708);
PE P1709(out_s1645, out_e1708, clk, rst, out_s1709, out_e1709, result1709);
PE P1710(out_s1646, out_e1709, clk, rst, out_s1710, out_e1710, result1710);
PE P1711(out_s1647, out_e1710, clk, rst, out_s1711, out_e1711, result1711);
PE P1712(out_s1648, out_e1711, clk, rst, out_s1712, out_e1712, result1712);
PE P1713(out_s1649, out_e1712, clk, rst, out_s1713, out_e1713, result1713);
PE P1714(out_s1650, out_e1713, clk, rst, out_s1714, out_e1714, result1714);
PE P1715(out_s1651, out_e1714, clk, rst, out_s1715, out_e1715, result1715);
PE P1716(out_s1652, out_e1715, clk, rst, out_s1716, out_e1716, result1716);
PE P1717(out_s1653, out_e1716, clk, rst, out_s1717, out_e1717, result1717);
PE P1718(out_s1654, out_e1717, clk, rst, out_s1718, out_e1718, result1718);
PE P1719(out_s1655, out_e1718, clk, rst, out_s1719, out_e1719, result1719);
PE P1720(out_s1656, out_e1719, clk, rst, out_s1720, out_e1720, result1720);
PE P1721(out_s1657, out_e1720, clk, rst, out_s1721, out_e1721, result1721);
PE P1722(out_s1658, out_e1721, clk, rst, out_s1722, out_e1722, result1722);
PE P1723(out_s1659, out_e1722, clk, rst, out_s1723, out_e1723, result1723);
PE P1724(out_s1660, out_e1723, clk, rst, out_s1724, out_e1724, result1724);
PE P1725(out_s1661, out_e1724, clk, rst, out_s1725, out_e1725, result1725);
PE P1726(out_s1662, out_e1725, clk, rst, out_s1726, out_e1726, result1726);
PE P1727(out_s1663, out_e1726, clk, rst, out_s1727, out_e1727, result1727);

PE P1729(out_s1665, out_e1728, clk, rst, out_s1729, out_e1729, result1729);
PE P1730(out_s1666, out_e1729, clk, rst, out_s1730, out_e1730, result1730);
PE P1731(out_s1667, out_e1730, clk, rst, out_s1731, out_e1731, result1731);
PE P1732(out_s1668, out_e1731, clk, rst, out_s1732, out_e1732, result1732);
PE P1733(out_s1669, out_e1732, clk, rst, out_s1733, out_e1733, result1733);
PE P1734(out_s1670, out_e1733, clk, rst, out_s1734, out_e1734, result1734);
PE P1735(out_s1671, out_e1734, clk, rst, out_s1735, out_e1735, result1735);
PE P1736(out_s1672, out_e1735, clk, rst, out_s1736, out_e1736, result1736);
PE P1737(out_s1673, out_e1736, clk, rst, out_s1737, out_e1737, result1737);
PE P1738(out_s1674, out_e1737, clk, rst, out_s1738, out_e1738, result1738);
PE P1739(out_s1675, out_e1738, clk, rst, out_s1739, out_e1739, result1739);
PE P1740(out_s1676, out_e1739, clk, rst, out_s1740, out_e1740, result1740);
PE P1741(out_s1677, out_e1740, clk, rst, out_s1741, out_e1741, result1741);
PE P1742(out_s1678, out_e1741, clk, rst, out_s1742, out_e1742, result1742);
PE P1743(out_s1679, out_e1742, clk, rst, out_s1743, out_e1743, result1743);
PE P1744(out_s1680, out_e1743, clk, rst, out_s1744, out_e1744, result1744);
PE P1745(out_s1681, out_e1744, clk, rst, out_s1745, out_e1745, result1745);
PE P1746(out_s1682, out_e1745, clk, rst, out_s1746, out_e1746, result1746);
PE P1747(out_s1683, out_e1746, clk, rst, out_s1747, out_e1747, result1747);
PE P1748(out_s1684, out_e1747, clk, rst, out_s1748, out_e1748, result1748);
PE P1749(out_s1685, out_e1748, clk, rst, out_s1749, out_e1749, result1749);
PE P1750(out_s1686, out_e1749, clk, rst, out_s1750, out_e1750, result1750);
PE P1751(out_s1687, out_e1750, clk, rst, out_s1751, out_e1751, result1751);
PE P1752(out_s1688, out_e1751, clk, rst, out_s1752, out_e1752, result1752);
PE P1753(out_s1689, out_e1752, clk, rst, out_s1753, out_e1753, result1753);
PE P1754(out_s1690, out_e1753, clk, rst, out_s1754, out_e1754, result1754);
PE P1755(out_s1691, out_e1754, clk, rst, out_s1755, out_e1755, result1755);
PE P1756(out_s1692, out_e1755, clk, rst, out_s1756, out_e1756, result1756);
PE P1757(out_s1693, out_e1756, clk, rst, out_s1757, out_e1757, result1757);
PE P1758(out_s1694, out_e1757, clk, rst, out_s1758, out_e1758, result1758);
PE P1759(out_s1695, out_e1758, clk, rst, out_s1759, out_e1759, result1759);
PE P1760(out_s1696, out_e1759, clk, rst, out_s1760, out_e1760, result1760);
PE P1761(out_s1697, out_e1760, clk, rst, out_s1761, out_e1761, result1761);
PE P1762(out_s1698, out_e1761, clk, rst, out_s1762, out_e1762, result1762);
PE P1763(out_s1699, out_e1762, clk, rst, out_s1763, out_e1763, result1763);
PE P1764(out_s1700, out_e1763, clk, rst, out_s1764, out_e1764, result1764);
PE P1765(out_s1701, out_e1764, clk, rst, out_s1765, out_e1765, result1765);
PE P1766(out_s1702, out_e1765, clk, rst, out_s1766, out_e1766, result1766);
PE P1767(out_s1703, out_e1766, clk, rst, out_s1767, out_e1767, result1767);
PE P1768(out_s1704, out_e1767, clk, rst, out_s1768, out_e1768, result1768);
PE P1769(out_s1705, out_e1768, clk, rst, out_s1769, out_e1769, result1769);
PE P1770(out_s1706, out_e1769, clk, rst, out_s1770, out_e1770, result1770);
PE P1771(out_s1707, out_e1770, clk, rst, out_s1771, out_e1771, result1771);
PE P1772(out_s1708, out_e1771, clk, rst, out_s1772, out_e1772, result1772);
PE P1773(out_s1709, out_e1772, clk, rst, out_s1773, out_e1773, result1773);
PE P1774(out_s1710, out_e1773, clk, rst, out_s1774, out_e1774, result1774);
PE P1775(out_s1711, out_e1774, clk, rst, out_s1775, out_e1775, result1775);
PE P1776(out_s1712, out_e1775, clk, rst, out_s1776, out_e1776, result1776);
PE P1777(out_s1713, out_e1776, clk, rst, out_s1777, out_e1777, result1777);
PE P1778(out_s1714, out_e1777, clk, rst, out_s1778, out_e1778, result1778);
PE P1779(out_s1715, out_e1778, clk, rst, out_s1779, out_e1779, result1779);
PE P1780(out_s1716, out_e1779, clk, rst, out_s1780, out_e1780, result1780);
PE P1781(out_s1717, out_e1780, clk, rst, out_s1781, out_e1781, result1781);
PE P1782(out_s1718, out_e1781, clk, rst, out_s1782, out_e1782, result1782);
PE P1783(out_s1719, out_e1782, clk, rst, out_s1783, out_e1783, result1783);
PE P1784(out_s1720, out_e1783, clk, rst, out_s1784, out_e1784, result1784);
PE P1785(out_s1721, out_e1784, clk, rst, out_s1785, out_e1785, result1785);
PE P1786(out_s1722, out_e1785, clk, rst, out_s1786, out_e1786, result1786);
PE P1787(out_s1723, out_e1786, clk, rst, out_s1787, out_e1787, result1787);
PE P1788(out_s1724, out_e1787, clk, rst, out_s1788, out_e1788, result1788);
PE P1789(out_s1725, out_e1788, clk, rst, out_s1789, out_e1789, result1789);
PE P1790(out_s1726, out_e1789, clk, rst, out_s1790, out_e1790, result1790);
PE P1791(out_s1727, out_e1790, clk, rst, out_s1791, out_e1791, result1791);

PE P1793(out_s1729, out_e1792, clk, rst, out_s1793, out_e1793, result1793);
PE P1794(out_s1730, out_e1793, clk, rst, out_s1794, out_e1794, result1794);
PE P1795(out_s1731, out_e1794, clk, rst, out_s1795, out_e1795, result1795);
PE P1796(out_s1732, out_e1795, clk, rst, out_s1796, out_e1796, result1796);
PE P1797(out_s1733, out_e1796, clk, rst, out_s1797, out_e1797, result1797);
PE P1798(out_s1734, out_e1797, clk, rst, out_s1798, out_e1798, result1798);
PE P1799(out_s1735, out_e1798, clk, rst, out_s1799, out_e1799, result1799);
PE P1800(out_s1736, out_e1799, clk, rst, out_s1800, out_e1800, result1800);
PE P1801(out_s1737, out_e1800, clk, rst, out_s1801, out_e1801, result1801);
PE P1802(out_s1738, out_e1801, clk, rst, out_s1802, out_e1802, result1802);
PE P1803(out_s1739, out_e1802, clk, rst, out_s1803, out_e1803, result1803);
PE P1804(out_s1740, out_e1803, clk, rst, out_s1804, out_e1804, result1804);
PE P1805(out_s1741, out_e1804, clk, rst, out_s1805, out_e1805, result1805);
PE P1806(out_s1742, out_e1805, clk, rst, out_s1806, out_e1806, result1806);
PE P1807(out_s1743, out_e1806, clk, rst, out_s1807, out_e1807, result1807);
PE P1808(out_s1744, out_e1807, clk, rst, out_s1808, out_e1808, result1808);
PE P1809(out_s1745, out_e1808, clk, rst, out_s1809, out_e1809, result1809);
PE P1810(out_s1746, out_e1809, clk, rst, out_s1810, out_e1810, result1810);
PE P1811(out_s1747, out_e1810, clk, rst, out_s1811, out_e1811, result1811);
PE P1812(out_s1748, out_e1811, clk, rst, out_s1812, out_e1812, result1812);
PE P1813(out_s1749, out_e1812, clk, rst, out_s1813, out_e1813, result1813);
PE P1814(out_s1750, out_e1813, clk, rst, out_s1814, out_e1814, result1814);
PE P1815(out_s1751, out_e1814, clk, rst, out_s1815, out_e1815, result1815);
PE P1816(out_s1752, out_e1815, clk, rst, out_s1816, out_e1816, result1816);
PE P1817(out_s1753, out_e1816, clk, rst, out_s1817, out_e1817, result1817);
PE P1818(out_s1754, out_e1817, clk, rst, out_s1818, out_e1818, result1818);
PE P1819(out_s1755, out_e1818, clk, rst, out_s1819, out_e1819, result1819);
PE P1820(out_s1756, out_e1819, clk, rst, out_s1820, out_e1820, result1820);
PE P1821(out_s1757, out_e1820, clk, rst, out_s1821, out_e1821, result1821);
PE P1822(out_s1758, out_e1821, clk, rst, out_s1822, out_e1822, result1822);
PE P1823(out_s1759, out_e1822, clk, rst, out_s1823, out_e1823, result1823);
PE P1824(out_s1760, out_e1823, clk, rst, out_s1824, out_e1824, result1824);
PE P1825(out_s1761, out_e1824, clk, rst, out_s1825, out_e1825, result1825);
PE P1826(out_s1762, out_e1825, clk, rst, out_s1826, out_e1826, result1826);
PE P1827(out_s1763, out_e1826, clk, rst, out_s1827, out_e1827, result1827);
PE P1828(out_s1764, out_e1827, clk, rst, out_s1828, out_e1828, result1828);
PE P1829(out_s1765, out_e1828, clk, rst, out_s1829, out_e1829, result1829);
PE P1830(out_s1766, out_e1829, clk, rst, out_s1830, out_e1830, result1830);
PE P1831(out_s1767, out_e1830, clk, rst, out_s1831, out_e1831, result1831);
PE P1832(out_s1768, out_e1831, clk, rst, out_s1832, out_e1832, result1832);
PE P1833(out_s1769, out_e1832, clk, rst, out_s1833, out_e1833, result1833);
PE P1834(out_s1770, out_e1833, clk, rst, out_s1834, out_e1834, result1834);
PE P1835(out_s1771, out_e1834, clk, rst, out_s1835, out_e1835, result1835);
PE P1836(out_s1772, out_e1835, clk, rst, out_s1836, out_e1836, result1836);
PE P1837(out_s1773, out_e1836, clk, rst, out_s1837, out_e1837, result1837);
PE P1838(out_s1774, out_e1837, clk, rst, out_s1838, out_e1838, result1838);
PE P1839(out_s1775, out_e1838, clk, rst, out_s1839, out_e1839, result1839);
PE P1840(out_s1776, out_e1839, clk, rst, out_s1840, out_e1840, result1840);
PE P1841(out_s1777, out_e1840, clk, rst, out_s1841, out_e1841, result1841);
PE P1842(out_s1778, out_e1841, clk, rst, out_s1842, out_e1842, result1842);
PE P1843(out_s1779, out_e1842, clk, rst, out_s1843, out_e1843, result1843);
PE P1844(out_s1780, out_e1843, clk, rst, out_s1844, out_e1844, result1844);
PE P1845(out_s1781, out_e1844, clk, rst, out_s1845, out_e1845, result1845);
PE P1846(out_s1782, out_e1845, clk, rst, out_s1846, out_e1846, result1846);
PE P1847(out_s1783, out_e1846, clk, rst, out_s1847, out_e1847, result1847);
PE P1848(out_s1784, out_e1847, clk, rst, out_s1848, out_e1848, result1848);
PE P1849(out_s1785, out_e1848, clk, rst, out_s1849, out_e1849, result1849);
PE P1850(out_s1786, out_e1849, clk, rst, out_s1850, out_e1850, result1850);
PE P1851(out_s1787, out_e1850, clk, rst, out_s1851, out_e1851, result1851);
PE P1852(out_s1788, out_e1851, clk, rst, out_s1852, out_e1852, result1852);
PE P1853(out_s1789, out_e1852, clk, rst, out_s1853, out_e1853, result1853);
PE P1854(out_s1790, out_e1853, clk, rst, out_s1854, out_e1854, result1854);
PE P1855(out_s1791, out_e1854, clk, rst, out_s1855, out_e1855, result1855);

PE P1857(out_s1793, out_e1856, clk, rst, out_s1857, out_e1857, result1857);
PE P1858(out_s1794, out_e1857, clk, rst, out_s1858, out_e1858, result1858);
PE P1859(out_s1795, out_e1858, clk, rst, out_s1859, out_e1859, result1859);
PE P1860(out_s1796, out_e1859, clk, rst, out_s1860, out_e1860, result1860);
PE P1861(out_s1797, out_e1860, clk, rst, out_s1861, out_e1861, result1861);
PE P1862(out_s1798, out_e1861, clk, rst, out_s1862, out_e1862, result1862);
PE P1863(out_s1799, out_e1862, clk, rst, out_s1863, out_e1863, result1863);
PE P1864(out_s1800, out_e1863, clk, rst, out_s1864, out_e1864, result1864);
PE P1865(out_s1801, out_e1864, clk, rst, out_s1865, out_e1865, result1865);
PE P1866(out_s1802, out_e1865, clk, rst, out_s1866, out_e1866, result1866);
PE P1867(out_s1803, out_e1866, clk, rst, out_s1867, out_e1867, result1867);
PE P1868(out_s1804, out_e1867, clk, rst, out_s1868, out_e1868, result1868);
PE P1869(out_s1805, out_e1868, clk, rst, out_s1869, out_e1869, result1869);
PE P1870(out_s1806, out_e1869, clk, rst, out_s1870, out_e1870, result1870);
PE P1871(out_s1807, out_e1870, clk, rst, out_s1871, out_e1871, result1871);
PE P1872(out_s1808, out_e1871, clk, rst, out_s1872, out_e1872, result1872);
PE P1873(out_s1809, out_e1872, clk, rst, out_s1873, out_e1873, result1873);
PE P1874(out_s1810, out_e1873, clk, rst, out_s1874, out_e1874, result1874);
PE P1875(out_s1811, out_e1874, clk, rst, out_s1875, out_e1875, result1875);
PE P1876(out_s1812, out_e1875, clk, rst, out_s1876, out_e1876, result1876);
PE P1877(out_s1813, out_e1876, clk, rst, out_s1877, out_e1877, result1877);
PE P1878(out_s1814, out_e1877, clk, rst, out_s1878, out_e1878, result1878);
PE P1879(out_s1815, out_e1878, clk, rst, out_s1879, out_e1879, result1879);
PE P1880(out_s1816, out_e1879, clk, rst, out_s1880, out_e1880, result1880);
PE P1881(out_s1817, out_e1880, clk, rst, out_s1881, out_e1881, result1881);
PE P1882(out_s1818, out_e1881, clk, rst, out_s1882, out_e1882, result1882);
PE P1883(out_s1819, out_e1882, clk, rst, out_s1883, out_e1883, result1883);
PE P1884(out_s1820, out_e1883, clk, rst, out_s1884, out_e1884, result1884);
PE P1885(out_s1821, out_e1884, clk, rst, out_s1885, out_e1885, result1885);
PE P1886(out_s1822, out_e1885, clk, rst, out_s1886, out_e1886, result1886);
PE P1887(out_s1823, out_e1886, clk, rst, out_s1887, out_e1887, result1887);
PE P1888(out_s1824, out_e1887, clk, rst, out_s1888, out_e1888, result1888);
PE P1889(out_s1825, out_e1888, clk, rst, out_s1889, out_e1889, result1889);
PE P1890(out_s1826, out_e1889, clk, rst, out_s1890, out_e1890, result1890);
PE P1891(out_s1827, out_e1890, clk, rst, out_s1891, out_e1891, result1891);
PE P1892(out_s1828, out_e1891, clk, rst, out_s1892, out_e1892, result1892);
PE P1893(out_s1829, out_e1892, clk, rst, out_s1893, out_e1893, result1893);
PE P1894(out_s1830, out_e1893, clk, rst, out_s1894, out_e1894, result1894);
PE P1895(out_s1831, out_e1894, clk, rst, out_s1895, out_e1895, result1895);
PE P1896(out_s1832, out_e1895, clk, rst, out_s1896, out_e1896, result1896);
PE P1897(out_s1833, out_e1896, clk, rst, out_s1897, out_e1897, result1897);
PE P1898(out_s1834, out_e1897, clk, rst, out_s1898, out_e1898, result1898);
PE P1899(out_s1835, out_e1898, clk, rst, out_s1899, out_e1899, result1899);
PE P1900(out_s1836, out_e1899, clk, rst, out_s1900, out_e1900, result1900);
PE P1901(out_s1837, out_e1900, clk, rst, out_s1901, out_e1901, result1901);
PE P1902(out_s1838, out_e1901, clk, rst, out_s1902, out_e1902, result1902);
PE P1903(out_s1839, out_e1902, clk, rst, out_s1903, out_e1903, result1903);
PE P1904(out_s1840, out_e1903, clk, rst, out_s1904, out_e1904, result1904);
PE P1905(out_s1841, out_e1904, clk, rst, out_s1905, out_e1905, result1905);
PE P1906(out_s1842, out_e1905, clk, rst, out_s1906, out_e1906, result1906);
PE P1907(out_s1843, out_e1906, clk, rst, out_s1907, out_e1907, result1907);
PE P1908(out_s1844, out_e1907, clk, rst, out_s1908, out_e1908, result1908);
PE P1909(out_s1845, out_e1908, clk, rst, out_s1909, out_e1909, result1909);
PE P1910(out_s1846, out_e1909, clk, rst, out_s1910, out_e1910, result1910);
PE P1911(out_s1847, out_e1910, clk, rst, out_s1911, out_e1911, result1911);
PE P1912(out_s1848, out_e1911, clk, rst, out_s1912, out_e1912, result1912);
PE P1913(out_s1849, out_e1912, clk, rst, out_s1913, out_e1913, result1913);
PE P1914(out_s1850, out_e1913, clk, rst, out_s1914, out_e1914, result1914);
PE P1915(out_s1851, out_e1914, clk, rst, out_s1915, out_e1915, result1915);
PE P1916(out_s1852, out_e1915, clk, rst, out_s1916, out_e1916, result1916);
PE P1917(out_s1853, out_e1916, clk, rst, out_s1917, out_e1917, result1917);
PE P1918(out_s1854, out_e1917, clk, rst, out_s1918, out_e1918, result1918);
PE P1919(out_s1855, out_e1918, clk, rst, out_s1919, out_e1919, result1919);

PE P1921(out_s1857, out_e1920, clk, rst, out_s1921, out_e1921, result1921);
PE P1922(out_s1858, out_e1921, clk, rst, out_s1922, out_e1922, result1922);
PE P1923(out_s1859, out_e1922, clk, rst, out_s1923, out_e1923, result1923);
PE P1924(out_s1860, out_e1923, clk, rst, out_s1924, out_e1924, result1924);
PE P1925(out_s1861, out_e1924, clk, rst, out_s1925, out_e1925, result1925);
PE P1926(out_s1862, out_e1925, clk, rst, out_s1926, out_e1926, result1926);
PE P1927(out_s1863, out_e1926, clk, rst, out_s1927, out_e1927, result1927);
PE P1928(out_s1864, out_e1927, clk, rst, out_s1928, out_e1928, result1928);
PE P1929(out_s1865, out_e1928, clk, rst, out_s1929, out_e1929, result1929);
PE P1930(out_s1866, out_e1929, clk, rst, out_s1930, out_e1930, result1930);
PE P1931(out_s1867, out_e1930, clk, rst, out_s1931, out_e1931, result1931);
PE P1932(out_s1868, out_e1931, clk, rst, out_s1932, out_e1932, result1932);
PE P1933(out_s1869, out_e1932, clk, rst, out_s1933, out_e1933, result1933);
PE P1934(out_s1870, out_e1933, clk, rst, out_s1934, out_e1934, result1934);
PE P1935(out_s1871, out_e1934, clk, rst, out_s1935, out_e1935, result1935);
PE P1936(out_s1872, out_e1935, clk, rst, out_s1936, out_e1936, result1936);
PE P1937(out_s1873, out_e1936, clk, rst, out_s1937, out_e1937, result1937);
PE P1938(out_s1874, out_e1937, clk, rst, out_s1938, out_e1938, result1938);
PE P1939(out_s1875, out_e1938, clk, rst, out_s1939, out_e1939, result1939);
PE P1940(out_s1876, out_e1939, clk, rst, out_s1940, out_e1940, result1940);
PE P1941(out_s1877, out_e1940, clk, rst, out_s1941, out_e1941, result1941);
PE P1942(out_s1878, out_e1941, clk, rst, out_s1942, out_e1942, result1942);
PE P1943(out_s1879, out_e1942, clk, rst, out_s1943, out_e1943, result1943);
PE P1944(out_s1880, out_e1943, clk, rst, out_s1944, out_e1944, result1944);
PE P1945(out_s1881, out_e1944, clk, rst, out_s1945, out_e1945, result1945);
PE P1946(out_s1882, out_e1945, clk, rst, out_s1946, out_e1946, result1946);
PE P1947(out_s1883, out_e1946, clk, rst, out_s1947, out_e1947, result1947);
PE P1948(out_s1884, out_e1947, clk, rst, out_s1948, out_e1948, result1948);
PE P1949(out_s1885, out_e1948, clk, rst, out_s1949, out_e1949, result1949);
PE P1950(out_s1886, out_e1949, clk, rst, out_s1950, out_e1950, result1950);
PE P1951(out_s1887, out_e1950, clk, rst, out_s1951, out_e1951, result1951);
PE P1952(out_s1888, out_e1951, clk, rst, out_s1952, out_e1952, result1952);
PE P1953(out_s1889, out_e1952, clk, rst, out_s1953, out_e1953, result1953);
PE P1954(out_s1890, out_e1953, clk, rst, out_s1954, out_e1954, result1954);
PE P1955(out_s1891, out_e1954, clk, rst, out_s1955, out_e1955, result1955);
PE P1956(out_s1892, out_e1955, clk, rst, out_s1956, out_e1956, result1956);
PE P1957(out_s1893, out_e1956, clk, rst, out_s1957, out_e1957, result1957);
PE P1958(out_s1894, out_e1957, clk, rst, out_s1958, out_e1958, result1958);
PE P1959(out_s1895, out_e1958, clk, rst, out_s1959, out_e1959, result1959);
PE P1960(out_s1896, out_e1959, clk, rst, out_s1960, out_e1960, result1960);
PE P1961(out_s1897, out_e1960, clk, rst, out_s1961, out_e1961, result1961);
PE P1962(out_s1898, out_e1961, clk, rst, out_s1962, out_e1962, result1962);
PE P1963(out_s1899, out_e1962, clk, rst, out_s1963, out_e1963, result1963);
PE P1964(out_s1900, out_e1963, clk, rst, out_s1964, out_e1964, result1964);
PE P1965(out_s1901, out_e1964, clk, rst, out_s1965, out_e1965, result1965);
PE P1966(out_s1902, out_e1965, clk, rst, out_s1966, out_e1966, result1966);
PE P1967(out_s1903, out_e1966, clk, rst, out_s1967, out_e1967, result1967);
PE P1968(out_s1904, out_e1967, clk, rst, out_s1968, out_e1968, result1968);
PE P1969(out_s1905, out_e1968, clk, rst, out_s1969, out_e1969, result1969);
PE P1970(out_s1906, out_e1969, clk, rst, out_s1970, out_e1970, result1970);
PE P1971(out_s1907, out_e1970, clk, rst, out_s1971, out_e1971, result1971);
PE P1972(out_s1908, out_e1971, clk, rst, out_s1972, out_e1972, result1972);
PE P1973(out_s1909, out_e1972, clk, rst, out_s1973, out_e1973, result1973);
PE P1974(out_s1910, out_e1973, clk, rst, out_s1974, out_e1974, result1974);
PE P1975(out_s1911, out_e1974, clk, rst, out_s1975, out_e1975, result1975);
PE P1976(out_s1912, out_e1975, clk, rst, out_s1976, out_e1976, result1976);
PE P1977(out_s1913, out_e1976, clk, rst, out_s1977, out_e1977, result1977);
PE P1978(out_s1914, out_e1977, clk, rst, out_s1978, out_e1978, result1978);
PE P1979(out_s1915, out_e1978, clk, rst, out_s1979, out_e1979, result1979);
PE P1980(out_s1916, out_e1979, clk, rst, out_s1980, out_e1980, result1980);
PE P1981(out_s1917, out_e1980, clk, rst, out_s1981, out_e1981, result1981);
PE P1982(out_s1918, out_e1981, clk, rst, out_s1982, out_e1982, result1982);
PE P1983(out_s1919, out_e1982, clk, rst, out_s1983, out_e1983, result1983);

PE P1985(out_s1921, out_e1984, clk, rst, out_s1985, out_e1985, result1985);
PE P1986(out_s1922, out_e1985, clk, rst, out_s1986, out_e1986, result1986);
PE P1987(out_s1923, out_e1986, clk, rst, out_s1987, out_e1987, result1987);
PE P1988(out_s1924, out_e1987, clk, rst, out_s1988, out_e1988, result1988);
PE P1989(out_s1925, out_e1988, clk, rst, out_s1989, out_e1989, result1989);
PE P1990(out_s1926, out_e1989, clk, rst, out_s1990, out_e1990, result1990);
PE P1991(out_s1927, out_e1990, clk, rst, out_s1991, out_e1991, result1991);
PE P1992(out_s1928, out_e1991, clk, rst, out_s1992, out_e1992, result1992);
PE P1993(out_s1929, out_e1992, clk, rst, out_s1993, out_e1993, result1993);
PE P1994(out_s1930, out_e1993, clk, rst, out_s1994, out_e1994, result1994);
PE P1995(out_s1931, out_e1994, clk, rst, out_s1995, out_e1995, result1995);
PE P1996(out_s1932, out_e1995, clk, rst, out_s1996, out_e1996, result1996);
PE P1997(out_s1933, out_e1996, clk, rst, out_s1997, out_e1997, result1997);
PE P1998(out_s1934, out_e1997, clk, rst, out_s1998, out_e1998, result1998);
PE P1999(out_s1935, out_e1998, clk, rst, out_s1999, out_e1999, result1999);
PE P2000(out_s1936, out_e1999, clk, rst, out_s2000, out_e2000, result2000);
PE P2001(out_s1937, out_e2000, clk, rst, out_s2001, out_e2001, result2001);
PE P2002(out_s1938, out_e2001, clk, rst, out_s2002, out_e2002, result2002);
PE P2003(out_s1939, out_e2002, clk, rst, out_s2003, out_e2003, result2003);
PE P2004(out_s1940, out_e2003, clk, rst, out_s2004, out_e2004, result2004);
PE P2005(out_s1941, out_e2004, clk, rst, out_s2005, out_e2005, result2005);
PE P2006(out_s1942, out_e2005, clk, rst, out_s2006, out_e2006, result2006);
PE P2007(out_s1943, out_e2006, clk, rst, out_s2007, out_e2007, result2007);
PE P2008(out_s1944, out_e2007, clk, rst, out_s2008, out_e2008, result2008);
PE P2009(out_s1945, out_e2008, clk, rst, out_s2009, out_e2009, result2009);
PE P2010(out_s1946, out_e2009, clk, rst, out_s2010, out_e2010, result2010);
PE P2011(out_s1947, out_e2010, clk, rst, out_s2011, out_e2011, result2011);
PE P2012(out_s1948, out_e2011, clk, rst, out_s2012, out_e2012, result2012);
PE P2013(out_s1949, out_e2012, clk, rst, out_s2013, out_e2013, result2013);
PE P2014(out_s1950, out_e2013, clk, rst, out_s2014, out_e2014, result2014);
PE P2015(out_s1951, out_e2014, clk, rst, out_s2015, out_e2015, result2015);
PE P2016(out_s1952, out_e2015, clk, rst, out_s2016, out_e2016, result2016);
PE P2017(out_s1953, out_e2016, clk, rst, out_s2017, out_e2017, result2017);
PE P2018(out_s1954, out_e2017, clk, rst, out_s2018, out_e2018, result2018);
PE P2019(out_s1955, out_e2018, clk, rst, out_s2019, out_e2019, result2019);
PE P2020(out_s1956, out_e2019, clk, rst, out_s2020, out_e2020, result2020);
PE P2021(out_s1957, out_e2020, clk, rst, out_s2021, out_e2021, result2021);
PE P2022(out_s1958, out_e2021, clk, rst, out_s2022, out_e2022, result2022);
PE P2023(out_s1959, out_e2022, clk, rst, out_s2023, out_e2023, result2023);
PE P2024(out_s1960, out_e2023, clk, rst, out_s2024, out_e2024, result2024);
PE P2025(out_s1961, out_e2024, clk, rst, out_s2025, out_e2025, result2025);
PE P2026(out_s1962, out_e2025, clk, rst, out_s2026, out_e2026, result2026);
PE P2027(out_s1963, out_e2026, clk, rst, out_s2027, out_e2027, result2027);
PE P2028(out_s1964, out_e2027, clk, rst, out_s2028, out_e2028, result2028);
PE P2029(out_s1965, out_e2028, clk, rst, out_s2029, out_e2029, result2029);
PE P2030(out_s1966, out_e2029, clk, rst, out_s2030, out_e2030, result2030);
PE P2031(out_s1967, out_e2030, clk, rst, out_s2031, out_e2031, result2031);
PE P2032(out_s1968, out_e2031, clk, rst, out_s2032, out_e2032, result2032);
PE P2033(out_s1969, out_e2032, clk, rst, out_s2033, out_e2033, result2033);
PE P2034(out_s1970, out_e2033, clk, rst, out_s2034, out_e2034, result2034);
PE P2035(out_s1971, out_e2034, clk, rst, out_s2035, out_e2035, result2035);
PE P2036(out_s1972, out_e2035, clk, rst, out_s2036, out_e2036, result2036);
PE P2037(out_s1973, out_e2036, clk, rst, out_s2037, out_e2037, result2037);
PE P2038(out_s1974, out_e2037, clk, rst, out_s2038, out_e2038, result2038);
PE P2039(out_s1975, out_e2038, clk, rst, out_s2039, out_e2039, result2039);
PE P2040(out_s1976, out_e2039, clk, rst, out_s2040, out_e2040, result2040);
PE P2041(out_s1977, out_e2040, clk, rst, out_s2041, out_e2041, result2041);
PE P2042(out_s1978, out_e2041, clk, rst, out_s2042, out_e2042, result2042);
PE P2043(out_s1979, out_e2042, clk, rst, out_s2043, out_e2043, result2043);
PE P2044(out_s1980, out_e2043, clk, rst, out_s2044, out_e2044, result2044);
PE P2045(out_s1981, out_e2044, clk, rst, out_s2045, out_e2045, result2045);
PE P2046(out_s1982, out_e2045, clk, rst, out_s2046, out_e2046, result2046);
PE P2047(out_s1983, out_e2046, clk, rst, out_s2047, out_e2047, result2047);

PE P2049(out_s1985, out_e2048, clk, rst, out_s2049, out_e2049, result2049);
PE P2050(out_s1986, out_e2049, clk, rst, out_s2050, out_e2050, result2050);
PE P2051(out_s1987, out_e2050, clk, rst, out_s2051, out_e2051, result2051);
PE P2052(out_s1988, out_e2051, clk, rst, out_s2052, out_e2052, result2052);
PE P2053(out_s1989, out_e2052, clk, rst, out_s2053, out_e2053, result2053);
PE P2054(out_s1990, out_e2053, clk, rst, out_s2054, out_e2054, result2054);
PE P2055(out_s1991, out_e2054, clk, rst, out_s2055, out_e2055, result2055);
PE P2056(out_s1992, out_e2055, clk, rst, out_s2056, out_e2056, result2056);
PE P2057(out_s1993, out_e2056, clk, rst, out_s2057, out_e2057, result2057);
PE P2058(out_s1994, out_e2057, clk, rst, out_s2058, out_e2058, result2058);
PE P2059(out_s1995, out_e2058, clk, rst, out_s2059, out_e2059, result2059);
PE P2060(out_s1996, out_e2059, clk, rst, out_s2060, out_e2060, result2060);
PE P2061(out_s1997, out_e2060, clk, rst, out_s2061, out_e2061, result2061);
PE P2062(out_s1998, out_e2061, clk, rst, out_s2062, out_e2062, result2062);
PE P2063(out_s1999, out_e2062, clk, rst, out_s2063, out_e2063, result2063);
PE P2064(out_s2000, out_e2063, clk, rst, out_s2064, out_e2064, result2064);
PE P2065(out_s2001, out_e2064, clk, rst, out_s2065, out_e2065, result2065);
PE P2066(out_s2002, out_e2065, clk, rst, out_s2066, out_e2066, result2066);
PE P2067(out_s2003, out_e2066, clk, rst, out_s2067, out_e2067, result2067);
PE P2068(out_s2004, out_e2067, clk, rst, out_s2068, out_e2068, result2068);
PE P2069(out_s2005, out_e2068, clk, rst, out_s2069, out_e2069, result2069);
PE P2070(out_s2006, out_e2069, clk, rst, out_s2070, out_e2070, result2070);
PE P2071(out_s2007, out_e2070, clk, rst, out_s2071, out_e2071, result2071);
PE P2072(out_s2008, out_e2071, clk, rst, out_s2072, out_e2072, result2072);
PE P2073(out_s2009, out_e2072, clk, rst, out_s2073, out_e2073, result2073);
PE P2074(out_s2010, out_e2073, clk, rst, out_s2074, out_e2074, result2074);
PE P2075(out_s2011, out_e2074, clk, rst, out_s2075, out_e2075, result2075);
PE P2076(out_s2012, out_e2075, clk, rst, out_s2076, out_e2076, result2076);
PE P2077(out_s2013, out_e2076, clk, rst, out_s2077, out_e2077, result2077);
PE P2078(out_s2014, out_e2077, clk, rst, out_s2078, out_e2078, result2078);
PE P2079(out_s2015, out_e2078, clk, rst, out_s2079, out_e2079, result2079);
PE P2080(out_s2016, out_e2079, clk, rst, out_s2080, out_e2080, result2080);
PE P2081(out_s2017, out_e2080, clk, rst, out_s2081, out_e2081, result2081);
PE P2082(out_s2018, out_e2081, clk, rst, out_s2082, out_e2082, result2082);
PE P2083(out_s2019, out_e2082, clk, rst, out_s2083, out_e2083, result2083);
PE P2084(out_s2020, out_e2083, clk, rst, out_s2084, out_e2084, result2084);
PE P2085(out_s2021, out_e2084, clk, rst, out_s2085, out_e2085, result2085);
PE P2086(out_s2022, out_e2085, clk, rst, out_s2086, out_e2086, result2086);
PE P2087(out_s2023, out_e2086, clk, rst, out_s2087, out_e2087, result2087);
PE P2088(out_s2024, out_e2087, clk, rst, out_s2088, out_e2088, result2088);
PE P2089(out_s2025, out_e2088, clk, rst, out_s2089, out_e2089, result2089);
PE P2090(out_s2026, out_e2089, clk, rst, out_s2090, out_e2090, result2090);
PE P2091(out_s2027, out_e2090, clk, rst, out_s2091, out_e2091, result2091);
PE P2092(out_s2028, out_e2091, clk, rst, out_s2092, out_e2092, result2092);
PE P2093(out_s2029, out_e2092, clk, rst, out_s2093, out_e2093, result2093);
PE P2094(out_s2030, out_e2093, clk, rst, out_s2094, out_e2094, result2094);
PE P2095(out_s2031, out_e2094, clk, rst, out_s2095, out_e2095, result2095);
PE P2096(out_s2032, out_e2095, clk, rst, out_s2096, out_e2096, result2096);
PE P2097(out_s2033, out_e2096, clk, rst, out_s2097, out_e2097, result2097);
PE P2098(out_s2034, out_e2097, clk, rst, out_s2098, out_e2098, result2098);
PE P2099(out_s2035, out_e2098, clk, rst, out_s2099, out_e2099, result2099);
PE P2100(out_s2036, out_e2099, clk, rst, out_s2100, out_e2100, result2100);
PE P2101(out_s2037, out_e2100, clk, rst, out_s2101, out_e2101, result2101);
PE P2102(out_s2038, out_e2101, clk, rst, out_s2102, out_e2102, result2102);
PE P2103(out_s2039, out_e2102, clk, rst, out_s2103, out_e2103, result2103);
PE P2104(out_s2040, out_e2103, clk, rst, out_s2104, out_e2104, result2104);
PE P2105(out_s2041, out_e2104, clk, rst, out_s2105, out_e2105, result2105);
PE P2106(out_s2042, out_e2105, clk, rst, out_s2106, out_e2106, result2106);
PE P2107(out_s2043, out_e2106, clk, rst, out_s2107, out_e2107, result2107);
PE P2108(out_s2044, out_e2107, clk, rst, out_s2108, out_e2108, result2108);
PE P2109(out_s2045, out_e2108, clk, rst, out_s2109, out_e2109, result2109);
PE P2110(out_s2046, out_e2109, clk, rst, out_s2110, out_e2110, result2110);
PE P2111(out_s2047, out_e2110, clk, rst, out_s2111, out_e2111, result2111);

PE P2113(out_s2049, out_e2112, clk, rst, out_s2113, out_e2113, result2113);
PE P2114(out_s2050, out_e2113, clk, rst, out_s2114, out_e2114, result2114);
PE P2115(out_s2051, out_e2114, clk, rst, out_s2115, out_e2115, result2115);
PE P2116(out_s2052, out_e2115, clk, rst, out_s2116, out_e2116, result2116);
PE P2117(out_s2053, out_e2116, clk, rst, out_s2117, out_e2117, result2117);
PE P2118(out_s2054, out_e2117, clk, rst, out_s2118, out_e2118, result2118);
PE P2119(out_s2055, out_e2118, clk, rst, out_s2119, out_e2119, result2119);
PE P2120(out_s2056, out_e2119, clk, rst, out_s2120, out_e2120, result2120);
PE P2121(out_s2057, out_e2120, clk, rst, out_s2121, out_e2121, result2121);
PE P2122(out_s2058, out_e2121, clk, rst, out_s2122, out_e2122, result2122);
PE P2123(out_s2059, out_e2122, clk, rst, out_s2123, out_e2123, result2123);
PE P2124(out_s2060, out_e2123, clk, rst, out_s2124, out_e2124, result2124);
PE P2125(out_s2061, out_e2124, clk, rst, out_s2125, out_e2125, result2125);
PE P2126(out_s2062, out_e2125, clk, rst, out_s2126, out_e2126, result2126);
PE P2127(out_s2063, out_e2126, clk, rst, out_s2127, out_e2127, result2127);
PE P2128(out_s2064, out_e2127, clk, rst, out_s2128, out_e2128, result2128);
PE P2129(out_s2065, out_e2128, clk, rst, out_s2129, out_e2129, result2129);
PE P2130(out_s2066, out_e2129, clk, rst, out_s2130, out_e2130, result2130);
PE P2131(out_s2067, out_e2130, clk, rst, out_s2131, out_e2131, result2131);
PE P2132(out_s2068, out_e2131, clk, rst, out_s2132, out_e2132, result2132);
PE P2133(out_s2069, out_e2132, clk, rst, out_s2133, out_e2133, result2133);
PE P2134(out_s2070, out_e2133, clk, rst, out_s2134, out_e2134, result2134);
PE P2135(out_s2071, out_e2134, clk, rst, out_s2135, out_e2135, result2135);
PE P2136(out_s2072, out_e2135, clk, rst, out_s2136, out_e2136, result2136);
PE P2137(out_s2073, out_e2136, clk, rst, out_s2137, out_e2137, result2137);
PE P2138(out_s2074, out_e2137, clk, rst, out_s2138, out_e2138, result2138);
PE P2139(out_s2075, out_e2138, clk, rst, out_s2139, out_e2139, result2139);
PE P2140(out_s2076, out_e2139, clk, rst, out_s2140, out_e2140, result2140);
PE P2141(out_s2077, out_e2140, clk, rst, out_s2141, out_e2141, result2141);
PE P2142(out_s2078, out_e2141, clk, rst, out_s2142, out_e2142, result2142);
PE P2143(out_s2079, out_e2142, clk, rst, out_s2143, out_e2143, result2143);
PE P2144(out_s2080, out_e2143, clk, rst, out_s2144, out_e2144, result2144);
PE P2145(out_s2081, out_e2144, clk, rst, out_s2145, out_e2145, result2145);
PE P2146(out_s2082, out_e2145, clk, rst, out_s2146, out_e2146, result2146);
PE P2147(out_s2083, out_e2146, clk, rst, out_s2147, out_e2147, result2147);
PE P2148(out_s2084, out_e2147, clk, rst, out_s2148, out_e2148, result2148);
PE P2149(out_s2085, out_e2148, clk, rst, out_s2149, out_e2149, result2149);
PE P2150(out_s2086, out_e2149, clk, rst, out_s2150, out_e2150, result2150);
PE P2151(out_s2087, out_e2150, clk, rst, out_s2151, out_e2151, result2151);
PE P2152(out_s2088, out_e2151, clk, rst, out_s2152, out_e2152, result2152);
PE P2153(out_s2089, out_e2152, clk, rst, out_s2153, out_e2153, result2153);
PE P2154(out_s2090, out_e2153, clk, rst, out_s2154, out_e2154, result2154);
PE P2155(out_s2091, out_e2154, clk, rst, out_s2155, out_e2155, result2155);
PE P2156(out_s2092, out_e2155, clk, rst, out_s2156, out_e2156, result2156);
PE P2157(out_s2093, out_e2156, clk, rst, out_s2157, out_e2157, result2157);
PE P2158(out_s2094, out_e2157, clk, rst, out_s2158, out_e2158, result2158);
PE P2159(out_s2095, out_e2158, clk, rst, out_s2159, out_e2159, result2159);
PE P2160(out_s2096, out_e2159, clk, rst, out_s2160, out_e2160, result2160);
PE P2161(out_s2097, out_e2160, clk, rst, out_s2161, out_e2161, result2161);
PE P2162(out_s2098, out_e2161, clk, rst, out_s2162, out_e2162, result2162);
PE P2163(out_s2099, out_e2162, clk, rst, out_s2163, out_e2163, result2163);
PE P2164(out_s2100, out_e2163, clk, rst, out_s2164, out_e2164, result2164);
PE P2165(out_s2101, out_e2164, clk, rst, out_s2165, out_e2165, result2165);
PE P2166(out_s2102, out_e2165, clk, rst, out_s2166, out_e2166, result2166);
PE P2167(out_s2103, out_e2166, clk, rst, out_s2167, out_e2167, result2167);
PE P2168(out_s2104, out_e2167, clk, rst, out_s2168, out_e2168, result2168);
PE P2169(out_s2105, out_e2168, clk, rst, out_s2169, out_e2169, result2169);
PE P2170(out_s2106, out_e2169, clk, rst, out_s2170, out_e2170, result2170);
PE P2171(out_s2107, out_e2170, clk, rst, out_s2171, out_e2171, result2171);
PE P2172(out_s2108, out_e2171, clk, rst, out_s2172, out_e2172, result2172);
PE P2173(out_s2109, out_e2172, clk, rst, out_s2173, out_e2173, result2173);
PE P2174(out_s2110, out_e2173, clk, rst, out_s2174, out_e2174, result2174);
PE P2175(out_s2111, out_e2174, clk, rst, out_s2175, out_e2175, result2175);

PE P2177(out_s2113, out_e2176, clk, rst, out_s2177, out_e2177, result2177);
PE P2178(out_s2114, out_e2177, clk, rst, out_s2178, out_e2178, result2178);
PE P2179(out_s2115, out_e2178, clk, rst, out_s2179, out_e2179, result2179);
PE P2180(out_s2116, out_e2179, clk, rst, out_s2180, out_e2180, result2180);
PE P2181(out_s2117, out_e2180, clk, rst, out_s2181, out_e2181, result2181);
PE P2182(out_s2118, out_e2181, clk, rst, out_s2182, out_e2182, result2182);
PE P2183(out_s2119, out_e2182, clk, rst, out_s2183, out_e2183, result2183);
PE P2184(out_s2120, out_e2183, clk, rst, out_s2184, out_e2184, result2184);
PE P2185(out_s2121, out_e2184, clk, rst, out_s2185, out_e2185, result2185);
PE P2186(out_s2122, out_e2185, clk, rst, out_s2186, out_e2186, result2186);
PE P2187(out_s2123, out_e2186, clk, rst, out_s2187, out_e2187, result2187);
PE P2188(out_s2124, out_e2187, clk, rst, out_s2188, out_e2188, result2188);
PE P2189(out_s2125, out_e2188, clk, rst, out_s2189, out_e2189, result2189);
PE P2190(out_s2126, out_e2189, clk, rst, out_s2190, out_e2190, result2190);
PE P2191(out_s2127, out_e2190, clk, rst, out_s2191, out_e2191, result2191);
PE P2192(out_s2128, out_e2191, clk, rst, out_s2192, out_e2192, result2192);
PE P2193(out_s2129, out_e2192, clk, rst, out_s2193, out_e2193, result2193);
PE P2194(out_s2130, out_e2193, clk, rst, out_s2194, out_e2194, result2194);
PE P2195(out_s2131, out_e2194, clk, rst, out_s2195, out_e2195, result2195);
PE P2196(out_s2132, out_e2195, clk, rst, out_s2196, out_e2196, result2196);
PE P2197(out_s2133, out_e2196, clk, rst, out_s2197, out_e2197, result2197);
PE P2198(out_s2134, out_e2197, clk, rst, out_s2198, out_e2198, result2198);
PE P2199(out_s2135, out_e2198, clk, rst, out_s2199, out_e2199, result2199);
PE P2200(out_s2136, out_e2199, clk, rst, out_s2200, out_e2200, result2200);
PE P2201(out_s2137, out_e2200, clk, rst, out_s2201, out_e2201, result2201);
PE P2202(out_s2138, out_e2201, clk, rst, out_s2202, out_e2202, result2202);
PE P2203(out_s2139, out_e2202, clk, rst, out_s2203, out_e2203, result2203);
PE P2204(out_s2140, out_e2203, clk, rst, out_s2204, out_e2204, result2204);
PE P2205(out_s2141, out_e2204, clk, rst, out_s2205, out_e2205, result2205);
PE P2206(out_s2142, out_e2205, clk, rst, out_s2206, out_e2206, result2206);
PE P2207(out_s2143, out_e2206, clk, rst, out_s2207, out_e2207, result2207);
PE P2208(out_s2144, out_e2207, clk, rst, out_s2208, out_e2208, result2208);
PE P2209(out_s2145, out_e2208, clk, rst, out_s2209, out_e2209, result2209);
PE P2210(out_s2146, out_e2209, clk, rst, out_s2210, out_e2210, result2210);
PE P2211(out_s2147, out_e2210, clk, rst, out_s2211, out_e2211, result2211);
PE P2212(out_s2148, out_e2211, clk, rst, out_s2212, out_e2212, result2212);
PE P2213(out_s2149, out_e2212, clk, rst, out_s2213, out_e2213, result2213);
PE P2214(out_s2150, out_e2213, clk, rst, out_s2214, out_e2214, result2214);
PE P2215(out_s2151, out_e2214, clk, rst, out_s2215, out_e2215, result2215);
PE P2216(out_s2152, out_e2215, clk, rst, out_s2216, out_e2216, result2216);
PE P2217(out_s2153, out_e2216, clk, rst, out_s2217, out_e2217, result2217);
PE P2218(out_s2154, out_e2217, clk, rst, out_s2218, out_e2218, result2218);
PE P2219(out_s2155, out_e2218, clk, rst, out_s2219, out_e2219, result2219);
PE P2220(out_s2156, out_e2219, clk, rst, out_s2220, out_e2220, result2220);
PE P2221(out_s2157, out_e2220, clk, rst, out_s2221, out_e2221, result2221);
PE P2222(out_s2158, out_e2221, clk, rst, out_s2222, out_e2222, result2222);
PE P2223(out_s2159, out_e2222, clk, rst, out_s2223, out_e2223, result2223);
PE P2224(out_s2160, out_e2223, clk, rst, out_s2224, out_e2224, result2224);
PE P2225(out_s2161, out_e2224, clk, rst, out_s2225, out_e2225, result2225);
PE P2226(out_s2162, out_e2225, clk, rst, out_s2226, out_e2226, result2226);
PE P2227(out_s2163, out_e2226, clk, rst, out_s2227, out_e2227, result2227);
PE P2228(out_s2164, out_e2227, clk, rst, out_s2228, out_e2228, result2228);
PE P2229(out_s2165, out_e2228, clk, rst, out_s2229, out_e2229, result2229);
PE P2230(out_s2166, out_e2229, clk, rst, out_s2230, out_e2230, result2230);
PE P2231(out_s2167, out_e2230, clk, rst, out_s2231, out_e2231, result2231);
PE P2232(out_s2168, out_e2231, clk, rst, out_s2232, out_e2232, result2232);
PE P2233(out_s2169, out_e2232, clk, rst, out_s2233, out_e2233, result2233);
PE P2234(out_s2170, out_e2233, clk, rst, out_s2234, out_e2234, result2234);
PE P2235(out_s2171, out_e2234, clk, rst, out_s2235, out_e2235, result2235);
PE P2236(out_s2172, out_e2235, clk, rst, out_s2236, out_e2236, result2236);
PE P2237(out_s2173, out_e2236, clk, rst, out_s2237, out_e2237, result2237);
PE P2238(out_s2174, out_e2237, clk, rst, out_s2238, out_e2238, result2238);
PE P2239(out_s2175, out_e2238, clk, rst, out_s2239, out_e2239, result2239);

PE P2241(out_s2177, out_e2240, clk, rst, out_s2241, out_e2241, result2241);
PE P2242(out_s2178, out_e2241, clk, rst, out_s2242, out_e2242, result2242);
PE P2243(out_s2179, out_e2242, clk, rst, out_s2243, out_e2243, result2243);
PE P2244(out_s2180, out_e2243, clk, rst, out_s2244, out_e2244, result2244);
PE P2245(out_s2181, out_e2244, clk, rst, out_s2245, out_e2245, result2245);
PE P2246(out_s2182, out_e2245, clk, rst, out_s2246, out_e2246, result2246);
PE P2247(out_s2183, out_e2246, clk, rst, out_s2247, out_e2247, result2247);
PE P2248(out_s2184, out_e2247, clk, rst, out_s2248, out_e2248, result2248);
PE P2249(out_s2185, out_e2248, clk, rst, out_s2249, out_e2249, result2249);
PE P2250(out_s2186, out_e2249, clk, rst, out_s2250, out_e2250, result2250);
PE P2251(out_s2187, out_e2250, clk, rst, out_s2251, out_e2251, result2251);
PE P2252(out_s2188, out_e2251, clk, rst, out_s2252, out_e2252, result2252);
PE P2253(out_s2189, out_e2252, clk, rst, out_s2253, out_e2253, result2253);
PE P2254(out_s2190, out_e2253, clk, rst, out_s2254, out_e2254, result2254);
PE P2255(out_s2191, out_e2254, clk, rst, out_s2255, out_e2255, result2255);
PE P2256(out_s2192, out_e2255, clk, rst, out_s2256, out_e2256, result2256);
PE P2257(out_s2193, out_e2256, clk, rst, out_s2257, out_e2257, result2257);
PE P2258(out_s2194, out_e2257, clk, rst, out_s2258, out_e2258, result2258);
PE P2259(out_s2195, out_e2258, clk, rst, out_s2259, out_e2259, result2259);
PE P2260(out_s2196, out_e2259, clk, rst, out_s2260, out_e2260, result2260);
PE P2261(out_s2197, out_e2260, clk, rst, out_s2261, out_e2261, result2261);
PE P2262(out_s2198, out_e2261, clk, rst, out_s2262, out_e2262, result2262);
PE P2263(out_s2199, out_e2262, clk, rst, out_s2263, out_e2263, result2263);
PE P2264(out_s2200, out_e2263, clk, rst, out_s2264, out_e2264, result2264);
PE P2265(out_s2201, out_e2264, clk, rst, out_s2265, out_e2265, result2265);
PE P2266(out_s2202, out_e2265, clk, rst, out_s2266, out_e2266, result2266);
PE P2267(out_s2203, out_e2266, clk, rst, out_s2267, out_e2267, result2267);
PE P2268(out_s2204, out_e2267, clk, rst, out_s2268, out_e2268, result2268);
PE P2269(out_s2205, out_e2268, clk, rst, out_s2269, out_e2269, result2269);
PE P2270(out_s2206, out_e2269, clk, rst, out_s2270, out_e2270, result2270);
PE P2271(out_s2207, out_e2270, clk, rst, out_s2271, out_e2271, result2271);
PE P2272(out_s2208, out_e2271, clk, rst, out_s2272, out_e2272, result2272);
PE P2273(out_s2209, out_e2272, clk, rst, out_s2273, out_e2273, result2273);
PE P2274(out_s2210, out_e2273, clk, rst, out_s2274, out_e2274, result2274);
PE P2275(out_s2211, out_e2274, clk, rst, out_s2275, out_e2275, result2275);
PE P2276(out_s2212, out_e2275, clk, rst, out_s2276, out_e2276, result2276);
PE P2277(out_s2213, out_e2276, clk, rst, out_s2277, out_e2277, result2277);
PE P2278(out_s2214, out_e2277, clk, rst, out_s2278, out_e2278, result2278);
PE P2279(out_s2215, out_e2278, clk, rst, out_s2279, out_e2279, result2279);
PE P2280(out_s2216, out_e2279, clk, rst, out_s2280, out_e2280, result2280);
PE P2281(out_s2217, out_e2280, clk, rst, out_s2281, out_e2281, result2281);
PE P2282(out_s2218, out_e2281, clk, rst, out_s2282, out_e2282, result2282);
PE P2283(out_s2219, out_e2282, clk, rst, out_s2283, out_e2283, result2283);
PE P2284(out_s2220, out_e2283, clk, rst, out_s2284, out_e2284, result2284);
PE P2285(out_s2221, out_e2284, clk, rst, out_s2285, out_e2285, result2285);
PE P2286(out_s2222, out_e2285, clk, rst, out_s2286, out_e2286, result2286);
PE P2287(out_s2223, out_e2286, clk, rst, out_s2287, out_e2287, result2287);
PE P2288(out_s2224, out_e2287, clk, rst, out_s2288, out_e2288, result2288);
PE P2289(out_s2225, out_e2288, clk, rst, out_s2289, out_e2289, result2289);
PE P2290(out_s2226, out_e2289, clk, rst, out_s2290, out_e2290, result2290);
PE P2291(out_s2227, out_e2290, clk, rst, out_s2291, out_e2291, result2291);
PE P2292(out_s2228, out_e2291, clk, rst, out_s2292, out_e2292, result2292);
PE P2293(out_s2229, out_e2292, clk, rst, out_s2293, out_e2293, result2293);
PE P2294(out_s2230, out_e2293, clk, rst, out_s2294, out_e2294, result2294);
PE P2295(out_s2231, out_e2294, clk, rst, out_s2295, out_e2295, result2295);
PE P2296(out_s2232, out_e2295, clk, rst, out_s2296, out_e2296, result2296);
PE P2297(out_s2233, out_e2296, clk, rst, out_s2297, out_e2297, result2297);
PE P2298(out_s2234, out_e2297, clk, rst, out_s2298, out_e2298, result2298);
PE P2299(out_s2235, out_e2298, clk, rst, out_s2299, out_e2299, result2299);
PE P2300(out_s2236, out_e2299, clk, rst, out_s2300, out_e2300, result2300);
PE P2301(out_s2237, out_e2300, clk, rst, out_s2301, out_e2301, result2301);
PE P2302(out_s2238, out_e2301, clk, rst, out_s2302, out_e2302, result2302);
PE P2303(out_s2239, out_e2302, clk, rst, out_s2303, out_e2303, result2303);

PE P2305(out_s2241, out_e2304, clk, rst, out_s2305, out_e2305, result2305);
PE P2306(out_s2242, out_e2305, clk, rst, out_s2306, out_e2306, result2306);
PE P2307(out_s2243, out_e2306, clk, rst, out_s2307, out_e2307, result2307);
PE P2308(out_s2244, out_e2307, clk, rst, out_s2308, out_e2308, result2308);
PE P2309(out_s2245, out_e2308, clk, rst, out_s2309, out_e2309, result2309);
PE P2310(out_s2246, out_e2309, clk, rst, out_s2310, out_e2310, result2310);
PE P2311(out_s2247, out_e2310, clk, rst, out_s2311, out_e2311, result2311);
PE P2312(out_s2248, out_e2311, clk, rst, out_s2312, out_e2312, result2312);
PE P2313(out_s2249, out_e2312, clk, rst, out_s2313, out_e2313, result2313);
PE P2314(out_s2250, out_e2313, clk, rst, out_s2314, out_e2314, result2314);
PE P2315(out_s2251, out_e2314, clk, rst, out_s2315, out_e2315, result2315);
PE P2316(out_s2252, out_e2315, clk, rst, out_s2316, out_e2316, result2316);
PE P2317(out_s2253, out_e2316, clk, rst, out_s2317, out_e2317, result2317);
PE P2318(out_s2254, out_e2317, clk, rst, out_s2318, out_e2318, result2318);
PE P2319(out_s2255, out_e2318, clk, rst, out_s2319, out_e2319, result2319);
PE P2320(out_s2256, out_e2319, clk, rst, out_s2320, out_e2320, result2320);
PE P2321(out_s2257, out_e2320, clk, rst, out_s2321, out_e2321, result2321);
PE P2322(out_s2258, out_e2321, clk, rst, out_s2322, out_e2322, result2322);
PE P2323(out_s2259, out_e2322, clk, rst, out_s2323, out_e2323, result2323);
PE P2324(out_s2260, out_e2323, clk, rst, out_s2324, out_e2324, result2324);
PE P2325(out_s2261, out_e2324, clk, rst, out_s2325, out_e2325, result2325);
PE P2326(out_s2262, out_e2325, clk, rst, out_s2326, out_e2326, result2326);
PE P2327(out_s2263, out_e2326, clk, rst, out_s2327, out_e2327, result2327);
PE P2328(out_s2264, out_e2327, clk, rst, out_s2328, out_e2328, result2328);
PE P2329(out_s2265, out_e2328, clk, rst, out_s2329, out_e2329, result2329);
PE P2330(out_s2266, out_e2329, clk, rst, out_s2330, out_e2330, result2330);
PE P2331(out_s2267, out_e2330, clk, rst, out_s2331, out_e2331, result2331);
PE P2332(out_s2268, out_e2331, clk, rst, out_s2332, out_e2332, result2332);
PE P2333(out_s2269, out_e2332, clk, rst, out_s2333, out_e2333, result2333);
PE P2334(out_s2270, out_e2333, clk, rst, out_s2334, out_e2334, result2334);
PE P2335(out_s2271, out_e2334, clk, rst, out_s2335, out_e2335, result2335);
PE P2336(out_s2272, out_e2335, clk, rst, out_s2336, out_e2336, result2336);
PE P2337(out_s2273, out_e2336, clk, rst, out_s2337, out_e2337, result2337);
PE P2338(out_s2274, out_e2337, clk, rst, out_s2338, out_e2338, result2338);
PE P2339(out_s2275, out_e2338, clk, rst, out_s2339, out_e2339, result2339);
PE P2340(out_s2276, out_e2339, clk, rst, out_s2340, out_e2340, result2340);
PE P2341(out_s2277, out_e2340, clk, rst, out_s2341, out_e2341, result2341);
PE P2342(out_s2278, out_e2341, clk, rst, out_s2342, out_e2342, result2342);
PE P2343(out_s2279, out_e2342, clk, rst, out_s2343, out_e2343, result2343);
PE P2344(out_s2280, out_e2343, clk, rst, out_s2344, out_e2344, result2344);
PE P2345(out_s2281, out_e2344, clk, rst, out_s2345, out_e2345, result2345);
PE P2346(out_s2282, out_e2345, clk, rst, out_s2346, out_e2346, result2346);
PE P2347(out_s2283, out_e2346, clk, rst, out_s2347, out_e2347, result2347);
PE P2348(out_s2284, out_e2347, clk, rst, out_s2348, out_e2348, result2348);
PE P2349(out_s2285, out_e2348, clk, rst, out_s2349, out_e2349, result2349);
PE P2350(out_s2286, out_e2349, clk, rst, out_s2350, out_e2350, result2350);
PE P2351(out_s2287, out_e2350, clk, rst, out_s2351, out_e2351, result2351);
PE P2352(out_s2288, out_e2351, clk, rst, out_s2352, out_e2352, result2352);
PE P2353(out_s2289, out_e2352, clk, rst, out_s2353, out_e2353, result2353);
PE P2354(out_s2290, out_e2353, clk, rst, out_s2354, out_e2354, result2354);
PE P2355(out_s2291, out_e2354, clk, rst, out_s2355, out_e2355, result2355);
PE P2356(out_s2292, out_e2355, clk, rst, out_s2356, out_e2356, result2356);
PE P2357(out_s2293, out_e2356, clk, rst, out_s2357, out_e2357, result2357);
PE P2358(out_s2294, out_e2357, clk, rst, out_s2358, out_e2358, result2358);
PE P2359(out_s2295, out_e2358, clk, rst, out_s2359, out_e2359, result2359);
PE P2360(out_s2296, out_e2359, clk, rst, out_s2360, out_e2360, result2360);
PE P2361(out_s2297, out_e2360, clk, rst, out_s2361, out_e2361, result2361);
PE P2362(out_s2298, out_e2361, clk, rst, out_s2362, out_e2362, result2362);
PE P2363(out_s2299, out_e2362, clk, rst, out_s2363, out_e2363, result2363);
PE P2364(out_s2300, out_e2363, clk, rst, out_s2364, out_e2364, result2364);
PE P2365(out_s2301, out_e2364, clk, rst, out_s2365, out_e2365, result2365);
PE P2366(out_s2302, out_e2365, clk, rst, out_s2366, out_e2366, result2366);
PE P2367(out_s2303, out_e2366, clk, rst, out_s2367, out_e2367, result2367);

PE P2369(out_s2305, out_e2368, clk, rst, out_s2369, out_e2369, result2369);
PE P2370(out_s2306, out_e2369, clk, rst, out_s2370, out_e2370, result2370);
PE P2371(out_s2307, out_e2370, clk, rst, out_s2371, out_e2371, result2371);
PE P2372(out_s2308, out_e2371, clk, rst, out_s2372, out_e2372, result2372);
PE P2373(out_s2309, out_e2372, clk, rst, out_s2373, out_e2373, result2373);
PE P2374(out_s2310, out_e2373, clk, rst, out_s2374, out_e2374, result2374);
PE P2375(out_s2311, out_e2374, clk, rst, out_s2375, out_e2375, result2375);
PE P2376(out_s2312, out_e2375, clk, rst, out_s2376, out_e2376, result2376);
PE P2377(out_s2313, out_e2376, clk, rst, out_s2377, out_e2377, result2377);
PE P2378(out_s2314, out_e2377, clk, rst, out_s2378, out_e2378, result2378);
PE P2379(out_s2315, out_e2378, clk, rst, out_s2379, out_e2379, result2379);
PE P2380(out_s2316, out_e2379, clk, rst, out_s2380, out_e2380, result2380);
PE P2381(out_s2317, out_e2380, clk, rst, out_s2381, out_e2381, result2381);
PE P2382(out_s2318, out_e2381, clk, rst, out_s2382, out_e2382, result2382);
PE P2383(out_s2319, out_e2382, clk, rst, out_s2383, out_e2383, result2383);
PE P2384(out_s2320, out_e2383, clk, rst, out_s2384, out_e2384, result2384);
PE P2385(out_s2321, out_e2384, clk, rst, out_s2385, out_e2385, result2385);
PE P2386(out_s2322, out_e2385, clk, rst, out_s2386, out_e2386, result2386);
PE P2387(out_s2323, out_e2386, clk, rst, out_s2387, out_e2387, result2387);
PE P2388(out_s2324, out_e2387, clk, rst, out_s2388, out_e2388, result2388);
PE P2389(out_s2325, out_e2388, clk, rst, out_s2389, out_e2389, result2389);
PE P2390(out_s2326, out_e2389, clk, rst, out_s2390, out_e2390, result2390);
PE P2391(out_s2327, out_e2390, clk, rst, out_s2391, out_e2391, result2391);
PE P2392(out_s2328, out_e2391, clk, rst, out_s2392, out_e2392, result2392);
PE P2393(out_s2329, out_e2392, clk, rst, out_s2393, out_e2393, result2393);
PE P2394(out_s2330, out_e2393, clk, rst, out_s2394, out_e2394, result2394);
PE P2395(out_s2331, out_e2394, clk, rst, out_s2395, out_e2395, result2395);
PE P2396(out_s2332, out_e2395, clk, rst, out_s2396, out_e2396, result2396);
PE P2397(out_s2333, out_e2396, clk, rst, out_s2397, out_e2397, result2397);
PE P2398(out_s2334, out_e2397, clk, rst, out_s2398, out_e2398, result2398);
PE P2399(out_s2335, out_e2398, clk, rst, out_s2399, out_e2399, result2399);
PE P2400(out_s2336, out_e2399, clk, rst, out_s2400, out_e2400, result2400);
PE P2401(out_s2337, out_e2400, clk, rst, out_s2401, out_e2401, result2401);
PE P2402(out_s2338, out_e2401, clk, rst, out_s2402, out_e2402, result2402);
PE P2403(out_s2339, out_e2402, clk, rst, out_s2403, out_e2403, result2403);
PE P2404(out_s2340, out_e2403, clk, rst, out_s2404, out_e2404, result2404);
PE P2405(out_s2341, out_e2404, clk, rst, out_s2405, out_e2405, result2405);
PE P2406(out_s2342, out_e2405, clk, rst, out_s2406, out_e2406, result2406);
PE P2407(out_s2343, out_e2406, clk, rst, out_s2407, out_e2407, result2407);
PE P2408(out_s2344, out_e2407, clk, rst, out_s2408, out_e2408, result2408);
PE P2409(out_s2345, out_e2408, clk, rst, out_s2409, out_e2409, result2409);
PE P2410(out_s2346, out_e2409, clk, rst, out_s2410, out_e2410, result2410);
PE P2411(out_s2347, out_e2410, clk, rst, out_s2411, out_e2411, result2411);
PE P2412(out_s2348, out_e2411, clk, rst, out_s2412, out_e2412, result2412);
PE P2413(out_s2349, out_e2412, clk, rst, out_s2413, out_e2413, result2413);
PE P2414(out_s2350, out_e2413, clk, rst, out_s2414, out_e2414, result2414);
PE P2415(out_s2351, out_e2414, clk, rst, out_s2415, out_e2415, result2415);
PE P2416(out_s2352, out_e2415, clk, rst, out_s2416, out_e2416, result2416);
PE P2417(out_s2353, out_e2416, clk, rst, out_s2417, out_e2417, result2417);
PE P2418(out_s2354, out_e2417, clk, rst, out_s2418, out_e2418, result2418);
PE P2419(out_s2355, out_e2418, clk, rst, out_s2419, out_e2419, result2419);
PE P2420(out_s2356, out_e2419, clk, rst, out_s2420, out_e2420, result2420);
PE P2421(out_s2357, out_e2420, clk, rst, out_s2421, out_e2421, result2421);
PE P2422(out_s2358, out_e2421, clk, rst, out_s2422, out_e2422, result2422);
PE P2423(out_s2359, out_e2422, clk, rst, out_s2423, out_e2423, result2423);
PE P2424(out_s2360, out_e2423, clk, rst, out_s2424, out_e2424, result2424);
PE P2425(out_s2361, out_e2424, clk, rst, out_s2425, out_e2425, result2425);
PE P2426(out_s2362, out_e2425, clk, rst, out_s2426, out_e2426, result2426);
PE P2427(out_s2363, out_e2426, clk, rst, out_s2427, out_e2427, result2427);
PE P2428(out_s2364, out_e2427, clk, rst, out_s2428, out_e2428, result2428);
PE P2429(out_s2365, out_e2428, clk, rst, out_s2429, out_e2429, result2429);
PE P2430(out_s2366, out_e2429, clk, rst, out_s2430, out_e2430, result2430);
PE P2431(out_s2367, out_e2430, clk, rst, out_s2431, out_e2431, result2431);

PE P2433(out_s2369, out_e2432, clk, rst, out_s2433, out_e2433, result2433);
PE P2434(out_s2370, out_e2433, clk, rst, out_s2434, out_e2434, result2434);
PE P2435(out_s2371, out_e2434, clk, rst, out_s2435, out_e2435, result2435);
PE P2436(out_s2372, out_e2435, clk, rst, out_s2436, out_e2436, result2436);
PE P2437(out_s2373, out_e2436, clk, rst, out_s2437, out_e2437, result2437);
PE P2438(out_s2374, out_e2437, clk, rst, out_s2438, out_e2438, result2438);
PE P2439(out_s2375, out_e2438, clk, rst, out_s2439, out_e2439, result2439);
PE P2440(out_s2376, out_e2439, clk, rst, out_s2440, out_e2440, result2440);
PE P2441(out_s2377, out_e2440, clk, rst, out_s2441, out_e2441, result2441);
PE P2442(out_s2378, out_e2441, clk, rst, out_s2442, out_e2442, result2442);
PE P2443(out_s2379, out_e2442, clk, rst, out_s2443, out_e2443, result2443);
PE P2444(out_s2380, out_e2443, clk, rst, out_s2444, out_e2444, result2444);
PE P2445(out_s2381, out_e2444, clk, rst, out_s2445, out_e2445, result2445);
PE P2446(out_s2382, out_e2445, clk, rst, out_s2446, out_e2446, result2446);
PE P2447(out_s2383, out_e2446, clk, rst, out_s2447, out_e2447, result2447);
PE P2448(out_s2384, out_e2447, clk, rst, out_s2448, out_e2448, result2448);
PE P2449(out_s2385, out_e2448, clk, rst, out_s2449, out_e2449, result2449);
PE P2450(out_s2386, out_e2449, clk, rst, out_s2450, out_e2450, result2450);
PE P2451(out_s2387, out_e2450, clk, rst, out_s2451, out_e2451, result2451);
PE P2452(out_s2388, out_e2451, clk, rst, out_s2452, out_e2452, result2452);
PE P2453(out_s2389, out_e2452, clk, rst, out_s2453, out_e2453, result2453);
PE P2454(out_s2390, out_e2453, clk, rst, out_s2454, out_e2454, result2454);
PE P2455(out_s2391, out_e2454, clk, rst, out_s2455, out_e2455, result2455);
PE P2456(out_s2392, out_e2455, clk, rst, out_s2456, out_e2456, result2456);
PE P2457(out_s2393, out_e2456, clk, rst, out_s2457, out_e2457, result2457);
PE P2458(out_s2394, out_e2457, clk, rst, out_s2458, out_e2458, result2458);
PE P2459(out_s2395, out_e2458, clk, rst, out_s2459, out_e2459, result2459);
PE P2460(out_s2396, out_e2459, clk, rst, out_s2460, out_e2460, result2460);
PE P2461(out_s2397, out_e2460, clk, rst, out_s2461, out_e2461, result2461);
PE P2462(out_s2398, out_e2461, clk, rst, out_s2462, out_e2462, result2462);
PE P2463(out_s2399, out_e2462, clk, rst, out_s2463, out_e2463, result2463);
PE P2464(out_s2400, out_e2463, clk, rst, out_s2464, out_e2464, result2464);
PE P2465(out_s2401, out_e2464, clk, rst, out_s2465, out_e2465, result2465);
PE P2466(out_s2402, out_e2465, clk, rst, out_s2466, out_e2466, result2466);
PE P2467(out_s2403, out_e2466, clk, rst, out_s2467, out_e2467, result2467);
PE P2468(out_s2404, out_e2467, clk, rst, out_s2468, out_e2468, result2468);
PE P2469(out_s2405, out_e2468, clk, rst, out_s2469, out_e2469, result2469);
PE P2470(out_s2406, out_e2469, clk, rst, out_s2470, out_e2470, result2470);
PE P2471(out_s2407, out_e2470, clk, rst, out_s2471, out_e2471, result2471);
PE P2472(out_s2408, out_e2471, clk, rst, out_s2472, out_e2472, result2472);
PE P2473(out_s2409, out_e2472, clk, rst, out_s2473, out_e2473, result2473);
PE P2474(out_s2410, out_e2473, clk, rst, out_s2474, out_e2474, result2474);
PE P2475(out_s2411, out_e2474, clk, rst, out_s2475, out_e2475, result2475);
PE P2476(out_s2412, out_e2475, clk, rst, out_s2476, out_e2476, result2476);
PE P2477(out_s2413, out_e2476, clk, rst, out_s2477, out_e2477, result2477);
PE P2478(out_s2414, out_e2477, clk, rst, out_s2478, out_e2478, result2478);
PE P2479(out_s2415, out_e2478, clk, rst, out_s2479, out_e2479, result2479);
PE P2480(out_s2416, out_e2479, clk, rst, out_s2480, out_e2480, result2480);
PE P2481(out_s2417, out_e2480, clk, rst, out_s2481, out_e2481, result2481);
PE P2482(out_s2418, out_e2481, clk, rst, out_s2482, out_e2482, result2482);
PE P2483(out_s2419, out_e2482, clk, rst, out_s2483, out_e2483, result2483);
PE P2484(out_s2420, out_e2483, clk, rst, out_s2484, out_e2484, result2484);
PE P2485(out_s2421, out_e2484, clk, rst, out_s2485, out_e2485, result2485);
PE P2486(out_s2422, out_e2485, clk, rst, out_s2486, out_e2486, result2486);
PE P2487(out_s2423, out_e2486, clk, rst, out_s2487, out_e2487, result2487);
PE P2488(out_s2424, out_e2487, clk, rst, out_s2488, out_e2488, result2488);
PE P2489(out_s2425, out_e2488, clk, rst, out_s2489, out_e2489, result2489);
PE P2490(out_s2426, out_e2489, clk, rst, out_s2490, out_e2490, result2490);
PE P2491(out_s2427, out_e2490, clk, rst, out_s2491, out_e2491, result2491);
PE P2492(out_s2428, out_e2491, clk, rst, out_s2492, out_e2492, result2492);
PE P2493(out_s2429, out_e2492, clk, rst, out_s2493, out_e2493, result2493);
PE P2494(out_s2430, out_e2493, clk, rst, out_s2494, out_e2494, result2494);
PE P2495(out_s2431, out_e2494, clk, rst, out_s2495, out_e2495, result2495);

PE P2497(out_s2433, out_e2496, clk, rst, out_s2497, out_e2497, result2497);
PE P2498(out_s2434, out_e2497, clk, rst, out_s2498, out_e2498, result2498);
PE P2499(out_s2435, out_e2498, clk, rst, out_s2499, out_e2499, result2499);
PE P2500(out_s2436, out_e2499, clk, rst, out_s2500, out_e2500, result2500);
PE P2501(out_s2437, out_e2500, clk, rst, out_s2501, out_e2501, result2501);
PE P2502(out_s2438, out_e2501, clk, rst, out_s2502, out_e2502, result2502);
PE P2503(out_s2439, out_e2502, clk, rst, out_s2503, out_e2503, result2503);
PE P2504(out_s2440, out_e2503, clk, rst, out_s2504, out_e2504, result2504);
PE P2505(out_s2441, out_e2504, clk, rst, out_s2505, out_e2505, result2505);
PE P2506(out_s2442, out_e2505, clk, rst, out_s2506, out_e2506, result2506);
PE P2507(out_s2443, out_e2506, clk, rst, out_s2507, out_e2507, result2507);
PE P2508(out_s2444, out_e2507, clk, rst, out_s2508, out_e2508, result2508);
PE P2509(out_s2445, out_e2508, clk, rst, out_s2509, out_e2509, result2509);
PE P2510(out_s2446, out_e2509, clk, rst, out_s2510, out_e2510, result2510);
PE P2511(out_s2447, out_e2510, clk, rst, out_s2511, out_e2511, result2511);
PE P2512(out_s2448, out_e2511, clk, rst, out_s2512, out_e2512, result2512);
PE P2513(out_s2449, out_e2512, clk, rst, out_s2513, out_e2513, result2513);
PE P2514(out_s2450, out_e2513, clk, rst, out_s2514, out_e2514, result2514);
PE P2515(out_s2451, out_e2514, clk, rst, out_s2515, out_e2515, result2515);
PE P2516(out_s2452, out_e2515, clk, rst, out_s2516, out_e2516, result2516);
PE P2517(out_s2453, out_e2516, clk, rst, out_s2517, out_e2517, result2517);
PE P2518(out_s2454, out_e2517, clk, rst, out_s2518, out_e2518, result2518);
PE P2519(out_s2455, out_e2518, clk, rst, out_s2519, out_e2519, result2519);
PE P2520(out_s2456, out_e2519, clk, rst, out_s2520, out_e2520, result2520);
PE P2521(out_s2457, out_e2520, clk, rst, out_s2521, out_e2521, result2521);
PE P2522(out_s2458, out_e2521, clk, rst, out_s2522, out_e2522, result2522);
PE P2523(out_s2459, out_e2522, clk, rst, out_s2523, out_e2523, result2523);
PE P2524(out_s2460, out_e2523, clk, rst, out_s2524, out_e2524, result2524);
PE P2525(out_s2461, out_e2524, clk, rst, out_s2525, out_e2525, result2525);
PE P2526(out_s2462, out_e2525, clk, rst, out_s2526, out_e2526, result2526);
PE P2527(out_s2463, out_e2526, clk, rst, out_s2527, out_e2527, result2527);
PE P2528(out_s2464, out_e2527, clk, rst, out_s2528, out_e2528, result2528);
PE P2529(out_s2465, out_e2528, clk, rst, out_s2529, out_e2529, result2529);
PE P2530(out_s2466, out_e2529, clk, rst, out_s2530, out_e2530, result2530);
PE P2531(out_s2467, out_e2530, clk, rst, out_s2531, out_e2531, result2531);
PE P2532(out_s2468, out_e2531, clk, rst, out_s2532, out_e2532, result2532);
PE P2533(out_s2469, out_e2532, clk, rst, out_s2533, out_e2533, result2533);
PE P2534(out_s2470, out_e2533, clk, rst, out_s2534, out_e2534, result2534);
PE P2535(out_s2471, out_e2534, clk, rst, out_s2535, out_e2535, result2535);
PE P2536(out_s2472, out_e2535, clk, rst, out_s2536, out_e2536, result2536);
PE P2537(out_s2473, out_e2536, clk, rst, out_s2537, out_e2537, result2537);
PE P2538(out_s2474, out_e2537, clk, rst, out_s2538, out_e2538, result2538);
PE P2539(out_s2475, out_e2538, clk, rst, out_s2539, out_e2539, result2539);
PE P2540(out_s2476, out_e2539, clk, rst, out_s2540, out_e2540, result2540);
PE P2541(out_s2477, out_e2540, clk, rst, out_s2541, out_e2541, result2541);
PE P2542(out_s2478, out_e2541, clk, rst, out_s2542, out_e2542, result2542);
PE P2543(out_s2479, out_e2542, clk, rst, out_s2543, out_e2543, result2543);
PE P2544(out_s2480, out_e2543, clk, rst, out_s2544, out_e2544, result2544);
PE P2545(out_s2481, out_e2544, clk, rst, out_s2545, out_e2545, result2545);
PE P2546(out_s2482, out_e2545, clk, rst, out_s2546, out_e2546, result2546);
PE P2547(out_s2483, out_e2546, clk, rst, out_s2547, out_e2547, result2547);
PE P2548(out_s2484, out_e2547, clk, rst, out_s2548, out_e2548, result2548);
PE P2549(out_s2485, out_e2548, clk, rst, out_s2549, out_e2549, result2549);
PE P2550(out_s2486, out_e2549, clk, rst, out_s2550, out_e2550, result2550);
PE P2551(out_s2487, out_e2550, clk, rst, out_s2551, out_e2551, result2551);
PE P2552(out_s2488, out_e2551, clk, rst, out_s2552, out_e2552, result2552);
PE P2553(out_s2489, out_e2552, clk, rst, out_s2553, out_e2553, result2553);
PE P2554(out_s2490, out_e2553, clk, rst, out_s2554, out_e2554, result2554);
PE P2555(out_s2491, out_e2554, clk, rst, out_s2555, out_e2555, result2555);
PE P2556(out_s2492, out_e2555, clk, rst, out_s2556, out_e2556, result2556);
PE P2557(out_s2493, out_e2556, clk, rst, out_s2557, out_e2557, result2557);
PE P2558(out_s2494, out_e2557, clk, rst, out_s2558, out_e2558, result2558);
PE P2559(out_s2495, out_e2558, clk, rst, out_s2559, out_e2559, result2559);

PE P2561(out_s2497, out_e2560, clk, rst, out_s2561, out_e2561, result2561);
PE P2562(out_s2498, out_e2561, clk, rst, out_s2562, out_e2562, result2562);
PE P2563(out_s2499, out_e2562, clk, rst, out_s2563, out_e2563, result2563);
PE P2564(out_s2500, out_e2563, clk, rst, out_s2564, out_e2564, result2564);
PE P2565(out_s2501, out_e2564, clk, rst, out_s2565, out_e2565, result2565);
PE P2566(out_s2502, out_e2565, clk, rst, out_s2566, out_e2566, result2566);
PE P2567(out_s2503, out_e2566, clk, rst, out_s2567, out_e2567, result2567);
PE P2568(out_s2504, out_e2567, clk, rst, out_s2568, out_e2568, result2568);
PE P2569(out_s2505, out_e2568, clk, rst, out_s2569, out_e2569, result2569);
PE P2570(out_s2506, out_e2569, clk, rst, out_s2570, out_e2570, result2570);
PE P2571(out_s2507, out_e2570, clk, rst, out_s2571, out_e2571, result2571);
PE P2572(out_s2508, out_e2571, clk, rst, out_s2572, out_e2572, result2572);
PE P2573(out_s2509, out_e2572, clk, rst, out_s2573, out_e2573, result2573);
PE P2574(out_s2510, out_e2573, clk, rst, out_s2574, out_e2574, result2574);
PE P2575(out_s2511, out_e2574, clk, rst, out_s2575, out_e2575, result2575);
PE P2576(out_s2512, out_e2575, clk, rst, out_s2576, out_e2576, result2576);
PE P2577(out_s2513, out_e2576, clk, rst, out_s2577, out_e2577, result2577);
PE P2578(out_s2514, out_e2577, clk, rst, out_s2578, out_e2578, result2578);
PE P2579(out_s2515, out_e2578, clk, rst, out_s2579, out_e2579, result2579);
PE P2580(out_s2516, out_e2579, clk, rst, out_s2580, out_e2580, result2580);
PE P2581(out_s2517, out_e2580, clk, rst, out_s2581, out_e2581, result2581);
PE P2582(out_s2518, out_e2581, clk, rst, out_s2582, out_e2582, result2582);
PE P2583(out_s2519, out_e2582, clk, rst, out_s2583, out_e2583, result2583);
PE P2584(out_s2520, out_e2583, clk, rst, out_s2584, out_e2584, result2584);
PE P2585(out_s2521, out_e2584, clk, rst, out_s2585, out_e2585, result2585);
PE P2586(out_s2522, out_e2585, clk, rst, out_s2586, out_e2586, result2586);
PE P2587(out_s2523, out_e2586, clk, rst, out_s2587, out_e2587, result2587);
PE P2588(out_s2524, out_e2587, clk, rst, out_s2588, out_e2588, result2588);
PE P2589(out_s2525, out_e2588, clk, rst, out_s2589, out_e2589, result2589);
PE P2590(out_s2526, out_e2589, clk, rst, out_s2590, out_e2590, result2590);
PE P2591(out_s2527, out_e2590, clk, rst, out_s2591, out_e2591, result2591);
PE P2592(out_s2528, out_e2591, clk, rst, out_s2592, out_e2592, result2592);
PE P2593(out_s2529, out_e2592, clk, rst, out_s2593, out_e2593, result2593);
PE P2594(out_s2530, out_e2593, clk, rst, out_s2594, out_e2594, result2594);
PE P2595(out_s2531, out_e2594, clk, rst, out_s2595, out_e2595, result2595);
PE P2596(out_s2532, out_e2595, clk, rst, out_s2596, out_e2596, result2596);
PE P2597(out_s2533, out_e2596, clk, rst, out_s2597, out_e2597, result2597);
PE P2598(out_s2534, out_e2597, clk, rst, out_s2598, out_e2598, result2598);
PE P2599(out_s2535, out_e2598, clk, rst, out_s2599, out_e2599, result2599);
PE P2600(out_s2536, out_e2599, clk, rst, out_s2600, out_e2600, result2600);
PE P2601(out_s2537, out_e2600, clk, rst, out_s2601, out_e2601, result2601);
PE P2602(out_s2538, out_e2601, clk, rst, out_s2602, out_e2602, result2602);
PE P2603(out_s2539, out_e2602, clk, rst, out_s2603, out_e2603, result2603);
PE P2604(out_s2540, out_e2603, clk, rst, out_s2604, out_e2604, result2604);
PE P2605(out_s2541, out_e2604, clk, rst, out_s2605, out_e2605, result2605);
PE P2606(out_s2542, out_e2605, clk, rst, out_s2606, out_e2606, result2606);
PE P2607(out_s2543, out_e2606, clk, rst, out_s2607, out_e2607, result2607);
PE P2608(out_s2544, out_e2607, clk, rst, out_s2608, out_e2608, result2608);
PE P2609(out_s2545, out_e2608, clk, rst, out_s2609, out_e2609, result2609);
PE P2610(out_s2546, out_e2609, clk, rst, out_s2610, out_e2610, result2610);
PE P2611(out_s2547, out_e2610, clk, rst, out_s2611, out_e2611, result2611);
PE P2612(out_s2548, out_e2611, clk, rst, out_s2612, out_e2612, result2612);
PE P2613(out_s2549, out_e2612, clk, rst, out_s2613, out_e2613, result2613);
PE P2614(out_s2550, out_e2613, clk, rst, out_s2614, out_e2614, result2614);
PE P2615(out_s2551, out_e2614, clk, rst, out_s2615, out_e2615, result2615);
PE P2616(out_s2552, out_e2615, clk, rst, out_s2616, out_e2616, result2616);
PE P2617(out_s2553, out_e2616, clk, rst, out_s2617, out_e2617, result2617);
PE P2618(out_s2554, out_e2617, clk, rst, out_s2618, out_e2618, result2618);
PE P2619(out_s2555, out_e2618, clk, rst, out_s2619, out_e2619, result2619);
PE P2620(out_s2556, out_e2619, clk, rst, out_s2620, out_e2620, result2620);
PE P2621(out_s2557, out_e2620, clk, rst, out_s2621, out_e2621, result2621);
PE P2622(out_s2558, out_e2621, clk, rst, out_s2622, out_e2622, result2622);
PE P2623(out_s2559, out_e2622, clk, rst, out_s2623, out_e2623, result2623);

PE P2625(out_s2561, out_e2624, clk, rst, out_s2625, out_e2625, result2625);
PE P2626(out_s2562, out_e2625, clk, rst, out_s2626, out_e2626, result2626);
PE P2627(out_s2563, out_e2626, clk, rst, out_s2627, out_e2627, result2627);
PE P2628(out_s2564, out_e2627, clk, rst, out_s2628, out_e2628, result2628);
PE P2629(out_s2565, out_e2628, clk, rst, out_s2629, out_e2629, result2629);
PE P2630(out_s2566, out_e2629, clk, rst, out_s2630, out_e2630, result2630);
PE P2631(out_s2567, out_e2630, clk, rst, out_s2631, out_e2631, result2631);
PE P2632(out_s2568, out_e2631, clk, rst, out_s2632, out_e2632, result2632);
PE P2633(out_s2569, out_e2632, clk, rst, out_s2633, out_e2633, result2633);
PE P2634(out_s2570, out_e2633, clk, rst, out_s2634, out_e2634, result2634);
PE P2635(out_s2571, out_e2634, clk, rst, out_s2635, out_e2635, result2635);
PE P2636(out_s2572, out_e2635, clk, rst, out_s2636, out_e2636, result2636);
PE P2637(out_s2573, out_e2636, clk, rst, out_s2637, out_e2637, result2637);
PE P2638(out_s2574, out_e2637, clk, rst, out_s2638, out_e2638, result2638);
PE P2639(out_s2575, out_e2638, clk, rst, out_s2639, out_e2639, result2639);
PE P2640(out_s2576, out_e2639, clk, rst, out_s2640, out_e2640, result2640);
PE P2641(out_s2577, out_e2640, clk, rst, out_s2641, out_e2641, result2641);
PE P2642(out_s2578, out_e2641, clk, rst, out_s2642, out_e2642, result2642);
PE P2643(out_s2579, out_e2642, clk, rst, out_s2643, out_e2643, result2643);
PE P2644(out_s2580, out_e2643, clk, rst, out_s2644, out_e2644, result2644);
PE P2645(out_s2581, out_e2644, clk, rst, out_s2645, out_e2645, result2645);
PE P2646(out_s2582, out_e2645, clk, rst, out_s2646, out_e2646, result2646);
PE P2647(out_s2583, out_e2646, clk, rst, out_s2647, out_e2647, result2647);
PE P2648(out_s2584, out_e2647, clk, rst, out_s2648, out_e2648, result2648);
PE P2649(out_s2585, out_e2648, clk, rst, out_s2649, out_e2649, result2649);
PE P2650(out_s2586, out_e2649, clk, rst, out_s2650, out_e2650, result2650);
PE P2651(out_s2587, out_e2650, clk, rst, out_s2651, out_e2651, result2651);
PE P2652(out_s2588, out_e2651, clk, rst, out_s2652, out_e2652, result2652);
PE P2653(out_s2589, out_e2652, clk, rst, out_s2653, out_e2653, result2653);
PE P2654(out_s2590, out_e2653, clk, rst, out_s2654, out_e2654, result2654);
PE P2655(out_s2591, out_e2654, clk, rst, out_s2655, out_e2655, result2655);
PE P2656(out_s2592, out_e2655, clk, rst, out_s2656, out_e2656, result2656);
PE P2657(out_s2593, out_e2656, clk, rst, out_s2657, out_e2657, result2657);
PE P2658(out_s2594, out_e2657, clk, rst, out_s2658, out_e2658, result2658);
PE P2659(out_s2595, out_e2658, clk, rst, out_s2659, out_e2659, result2659);
PE P2660(out_s2596, out_e2659, clk, rst, out_s2660, out_e2660, result2660);
PE P2661(out_s2597, out_e2660, clk, rst, out_s2661, out_e2661, result2661);
PE P2662(out_s2598, out_e2661, clk, rst, out_s2662, out_e2662, result2662);
PE P2663(out_s2599, out_e2662, clk, rst, out_s2663, out_e2663, result2663);
PE P2664(out_s2600, out_e2663, clk, rst, out_s2664, out_e2664, result2664);
PE P2665(out_s2601, out_e2664, clk, rst, out_s2665, out_e2665, result2665);
PE P2666(out_s2602, out_e2665, clk, rst, out_s2666, out_e2666, result2666);
PE P2667(out_s2603, out_e2666, clk, rst, out_s2667, out_e2667, result2667);
PE P2668(out_s2604, out_e2667, clk, rst, out_s2668, out_e2668, result2668);
PE P2669(out_s2605, out_e2668, clk, rst, out_s2669, out_e2669, result2669);
PE P2670(out_s2606, out_e2669, clk, rst, out_s2670, out_e2670, result2670);
PE P2671(out_s2607, out_e2670, clk, rst, out_s2671, out_e2671, result2671);
PE P2672(out_s2608, out_e2671, clk, rst, out_s2672, out_e2672, result2672);
PE P2673(out_s2609, out_e2672, clk, rst, out_s2673, out_e2673, result2673);
PE P2674(out_s2610, out_e2673, clk, rst, out_s2674, out_e2674, result2674);
PE P2675(out_s2611, out_e2674, clk, rst, out_s2675, out_e2675, result2675);
PE P2676(out_s2612, out_e2675, clk, rst, out_s2676, out_e2676, result2676);
PE P2677(out_s2613, out_e2676, clk, rst, out_s2677, out_e2677, result2677);
PE P2678(out_s2614, out_e2677, clk, rst, out_s2678, out_e2678, result2678);
PE P2679(out_s2615, out_e2678, clk, rst, out_s2679, out_e2679, result2679);
PE P2680(out_s2616, out_e2679, clk, rst, out_s2680, out_e2680, result2680);
PE P2681(out_s2617, out_e2680, clk, rst, out_s2681, out_e2681, result2681);
PE P2682(out_s2618, out_e2681, clk, rst, out_s2682, out_e2682, result2682);
PE P2683(out_s2619, out_e2682, clk, rst, out_s2683, out_e2683, result2683);
PE P2684(out_s2620, out_e2683, clk, rst, out_s2684, out_e2684, result2684);
PE P2685(out_s2621, out_e2684, clk, rst, out_s2685, out_e2685, result2685);
PE P2686(out_s2622, out_e2685, clk, rst, out_s2686, out_e2686, result2686);
PE P2687(out_s2623, out_e2686, clk, rst, out_s2687, out_e2687, result2687);

PE P2689(out_s2625, out_e2688, clk, rst, out_s2689, out_e2689, result2689);
PE P2690(out_s2626, out_e2689, clk, rst, out_s2690, out_e2690, result2690);
PE P2691(out_s2627, out_e2690, clk, rst, out_s2691, out_e2691, result2691);
PE P2692(out_s2628, out_e2691, clk, rst, out_s2692, out_e2692, result2692);
PE P2693(out_s2629, out_e2692, clk, rst, out_s2693, out_e2693, result2693);
PE P2694(out_s2630, out_e2693, clk, rst, out_s2694, out_e2694, result2694);
PE P2695(out_s2631, out_e2694, clk, rst, out_s2695, out_e2695, result2695);
PE P2696(out_s2632, out_e2695, clk, rst, out_s2696, out_e2696, result2696);
PE P2697(out_s2633, out_e2696, clk, rst, out_s2697, out_e2697, result2697);
PE P2698(out_s2634, out_e2697, clk, rst, out_s2698, out_e2698, result2698);
PE P2699(out_s2635, out_e2698, clk, rst, out_s2699, out_e2699, result2699);
PE P2700(out_s2636, out_e2699, clk, rst, out_s2700, out_e2700, result2700);
PE P2701(out_s2637, out_e2700, clk, rst, out_s2701, out_e2701, result2701);
PE P2702(out_s2638, out_e2701, clk, rst, out_s2702, out_e2702, result2702);
PE P2703(out_s2639, out_e2702, clk, rst, out_s2703, out_e2703, result2703);
PE P2704(out_s2640, out_e2703, clk, rst, out_s2704, out_e2704, result2704);
PE P2705(out_s2641, out_e2704, clk, rst, out_s2705, out_e2705, result2705);
PE P2706(out_s2642, out_e2705, clk, rst, out_s2706, out_e2706, result2706);
PE P2707(out_s2643, out_e2706, clk, rst, out_s2707, out_e2707, result2707);
PE P2708(out_s2644, out_e2707, clk, rst, out_s2708, out_e2708, result2708);
PE P2709(out_s2645, out_e2708, clk, rst, out_s2709, out_e2709, result2709);
PE P2710(out_s2646, out_e2709, clk, rst, out_s2710, out_e2710, result2710);
PE P2711(out_s2647, out_e2710, clk, rst, out_s2711, out_e2711, result2711);
PE P2712(out_s2648, out_e2711, clk, rst, out_s2712, out_e2712, result2712);
PE P2713(out_s2649, out_e2712, clk, rst, out_s2713, out_e2713, result2713);
PE P2714(out_s2650, out_e2713, clk, rst, out_s2714, out_e2714, result2714);
PE P2715(out_s2651, out_e2714, clk, rst, out_s2715, out_e2715, result2715);
PE P2716(out_s2652, out_e2715, clk, rst, out_s2716, out_e2716, result2716);
PE P2717(out_s2653, out_e2716, clk, rst, out_s2717, out_e2717, result2717);
PE P2718(out_s2654, out_e2717, clk, rst, out_s2718, out_e2718, result2718);
PE P2719(out_s2655, out_e2718, clk, rst, out_s2719, out_e2719, result2719);
PE P2720(out_s2656, out_e2719, clk, rst, out_s2720, out_e2720, result2720);
PE P2721(out_s2657, out_e2720, clk, rst, out_s2721, out_e2721, result2721);
PE P2722(out_s2658, out_e2721, clk, rst, out_s2722, out_e2722, result2722);
PE P2723(out_s2659, out_e2722, clk, rst, out_s2723, out_e2723, result2723);
PE P2724(out_s2660, out_e2723, clk, rst, out_s2724, out_e2724, result2724);
PE P2725(out_s2661, out_e2724, clk, rst, out_s2725, out_e2725, result2725);
PE P2726(out_s2662, out_e2725, clk, rst, out_s2726, out_e2726, result2726);
PE P2727(out_s2663, out_e2726, clk, rst, out_s2727, out_e2727, result2727);
PE P2728(out_s2664, out_e2727, clk, rst, out_s2728, out_e2728, result2728);
PE P2729(out_s2665, out_e2728, clk, rst, out_s2729, out_e2729, result2729);
PE P2730(out_s2666, out_e2729, clk, rst, out_s2730, out_e2730, result2730);
PE P2731(out_s2667, out_e2730, clk, rst, out_s2731, out_e2731, result2731);
PE P2732(out_s2668, out_e2731, clk, rst, out_s2732, out_e2732, result2732);
PE P2733(out_s2669, out_e2732, clk, rst, out_s2733, out_e2733, result2733);
PE P2734(out_s2670, out_e2733, clk, rst, out_s2734, out_e2734, result2734);
PE P2735(out_s2671, out_e2734, clk, rst, out_s2735, out_e2735, result2735);
PE P2736(out_s2672, out_e2735, clk, rst, out_s2736, out_e2736, result2736);
PE P2737(out_s2673, out_e2736, clk, rst, out_s2737, out_e2737, result2737);
PE P2738(out_s2674, out_e2737, clk, rst, out_s2738, out_e2738, result2738);
PE P2739(out_s2675, out_e2738, clk, rst, out_s2739, out_e2739, result2739);
PE P2740(out_s2676, out_e2739, clk, rst, out_s2740, out_e2740, result2740);
PE P2741(out_s2677, out_e2740, clk, rst, out_s2741, out_e2741, result2741);
PE P2742(out_s2678, out_e2741, clk, rst, out_s2742, out_e2742, result2742);
PE P2743(out_s2679, out_e2742, clk, rst, out_s2743, out_e2743, result2743);
PE P2744(out_s2680, out_e2743, clk, rst, out_s2744, out_e2744, result2744);
PE P2745(out_s2681, out_e2744, clk, rst, out_s2745, out_e2745, result2745);
PE P2746(out_s2682, out_e2745, clk, rst, out_s2746, out_e2746, result2746);
PE P2747(out_s2683, out_e2746, clk, rst, out_s2747, out_e2747, result2747);
PE P2748(out_s2684, out_e2747, clk, rst, out_s2748, out_e2748, result2748);
PE P2749(out_s2685, out_e2748, clk, rst, out_s2749, out_e2749, result2749);
PE P2750(out_s2686, out_e2749, clk, rst, out_s2750, out_e2750, result2750);
PE P2751(out_s2687, out_e2750, clk, rst, out_s2751, out_e2751, result2751);

PE P2753(out_s2689, out_e2752, clk, rst, out_s2753, out_e2753, result2753);
PE P2754(out_s2690, out_e2753, clk, rst, out_s2754, out_e2754, result2754);
PE P2755(out_s2691, out_e2754, clk, rst, out_s2755, out_e2755, result2755);
PE P2756(out_s2692, out_e2755, clk, rst, out_s2756, out_e2756, result2756);
PE P2757(out_s2693, out_e2756, clk, rst, out_s2757, out_e2757, result2757);
PE P2758(out_s2694, out_e2757, clk, rst, out_s2758, out_e2758, result2758);
PE P2759(out_s2695, out_e2758, clk, rst, out_s2759, out_e2759, result2759);
PE P2760(out_s2696, out_e2759, clk, rst, out_s2760, out_e2760, result2760);
PE P2761(out_s2697, out_e2760, clk, rst, out_s2761, out_e2761, result2761);
PE P2762(out_s2698, out_e2761, clk, rst, out_s2762, out_e2762, result2762);
PE P2763(out_s2699, out_e2762, clk, rst, out_s2763, out_e2763, result2763);
PE P2764(out_s2700, out_e2763, clk, rst, out_s2764, out_e2764, result2764);
PE P2765(out_s2701, out_e2764, clk, rst, out_s2765, out_e2765, result2765);
PE P2766(out_s2702, out_e2765, clk, rst, out_s2766, out_e2766, result2766);
PE P2767(out_s2703, out_e2766, clk, rst, out_s2767, out_e2767, result2767);
PE P2768(out_s2704, out_e2767, clk, rst, out_s2768, out_e2768, result2768);
PE P2769(out_s2705, out_e2768, clk, rst, out_s2769, out_e2769, result2769);
PE P2770(out_s2706, out_e2769, clk, rst, out_s2770, out_e2770, result2770);
PE P2771(out_s2707, out_e2770, clk, rst, out_s2771, out_e2771, result2771);
PE P2772(out_s2708, out_e2771, clk, rst, out_s2772, out_e2772, result2772);
PE P2773(out_s2709, out_e2772, clk, rst, out_s2773, out_e2773, result2773);
PE P2774(out_s2710, out_e2773, clk, rst, out_s2774, out_e2774, result2774);
PE P2775(out_s2711, out_e2774, clk, rst, out_s2775, out_e2775, result2775);
PE P2776(out_s2712, out_e2775, clk, rst, out_s2776, out_e2776, result2776);
PE P2777(out_s2713, out_e2776, clk, rst, out_s2777, out_e2777, result2777);
PE P2778(out_s2714, out_e2777, clk, rst, out_s2778, out_e2778, result2778);
PE P2779(out_s2715, out_e2778, clk, rst, out_s2779, out_e2779, result2779);
PE P2780(out_s2716, out_e2779, clk, rst, out_s2780, out_e2780, result2780);
PE P2781(out_s2717, out_e2780, clk, rst, out_s2781, out_e2781, result2781);
PE P2782(out_s2718, out_e2781, clk, rst, out_s2782, out_e2782, result2782);
PE P2783(out_s2719, out_e2782, clk, rst, out_s2783, out_e2783, result2783);
PE P2784(out_s2720, out_e2783, clk, rst, out_s2784, out_e2784, result2784);
PE P2785(out_s2721, out_e2784, clk, rst, out_s2785, out_e2785, result2785);
PE P2786(out_s2722, out_e2785, clk, rst, out_s2786, out_e2786, result2786);
PE P2787(out_s2723, out_e2786, clk, rst, out_s2787, out_e2787, result2787);
PE P2788(out_s2724, out_e2787, clk, rst, out_s2788, out_e2788, result2788);
PE P2789(out_s2725, out_e2788, clk, rst, out_s2789, out_e2789, result2789);
PE P2790(out_s2726, out_e2789, clk, rst, out_s2790, out_e2790, result2790);
PE P2791(out_s2727, out_e2790, clk, rst, out_s2791, out_e2791, result2791);
PE P2792(out_s2728, out_e2791, clk, rst, out_s2792, out_e2792, result2792);
PE P2793(out_s2729, out_e2792, clk, rst, out_s2793, out_e2793, result2793);
PE P2794(out_s2730, out_e2793, clk, rst, out_s2794, out_e2794, result2794);
PE P2795(out_s2731, out_e2794, clk, rst, out_s2795, out_e2795, result2795);
PE P2796(out_s2732, out_e2795, clk, rst, out_s2796, out_e2796, result2796);
PE P2797(out_s2733, out_e2796, clk, rst, out_s2797, out_e2797, result2797);
PE P2798(out_s2734, out_e2797, clk, rst, out_s2798, out_e2798, result2798);
PE P2799(out_s2735, out_e2798, clk, rst, out_s2799, out_e2799, result2799);
PE P2800(out_s2736, out_e2799, clk, rst, out_s2800, out_e2800, result2800);
PE P2801(out_s2737, out_e2800, clk, rst, out_s2801, out_e2801, result2801);
PE P2802(out_s2738, out_e2801, clk, rst, out_s2802, out_e2802, result2802);
PE P2803(out_s2739, out_e2802, clk, rst, out_s2803, out_e2803, result2803);
PE P2804(out_s2740, out_e2803, clk, rst, out_s2804, out_e2804, result2804);
PE P2805(out_s2741, out_e2804, clk, rst, out_s2805, out_e2805, result2805);
PE P2806(out_s2742, out_e2805, clk, rst, out_s2806, out_e2806, result2806);
PE P2807(out_s2743, out_e2806, clk, rst, out_s2807, out_e2807, result2807);
PE P2808(out_s2744, out_e2807, clk, rst, out_s2808, out_e2808, result2808);
PE P2809(out_s2745, out_e2808, clk, rst, out_s2809, out_e2809, result2809);
PE P2810(out_s2746, out_e2809, clk, rst, out_s2810, out_e2810, result2810);
PE P2811(out_s2747, out_e2810, clk, rst, out_s2811, out_e2811, result2811);
PE P2812(out_s2748, out_e2811, clk, rst, out_s2812, out_e2812, result2812);
PE P2813(out_s2749, out_e2812, clk, rst, out_s2813, out_e2813, result2813);
PE P2814(out_s2750, out_e2813, clk, rst, out_s2814, out_e2814, result2814);
PE P2815(out_s2751, out_e2814, clk, rst, out_s2815, out_e2815, result2815);

PE P2817(out_s2753, out_e2816, clk, rst, out_s2817, out_e2817, result2817);
PE P2818(out_s2754, out_e2817, clk, rst, out_s2818, out_e2818, result2818);
PE P2819(out_s2755, out_e2818, clk, rst, out_s2819, out_e2819, result2819);
PE P2820(out_s2756, out_e2819, clk, rst, out_s2820, out_e2820, result2820);
PE P2821(out_s2757, out_e2820, clk, rst, out_s2821, out_e2821, result2821);
PE P2822(out_s2758, out_e2821, clk, rst, out_s2822, out_e2822, result2822);
PE P2823(out_s2759, out_e2822, clk, rst, out_s2823, out_e2823, result2823);
PE P2824(out_s2760, out_e2823, clk, rst, out_s2824, out_e2824, result2824);
PE P2825(out_s2761, out_e2824, clk, rst, out_s2825, out_e2825, result2825);
PE P2826(out_s2762, out_e2825, clk, rst, out_s2826, out_e2826, result2826);
PE P2827(out_s2763, out_e2826, clk, rst, out_s2827, out_e2827, result2827);
PE P2828(out_s2764, out_e2827, clk, rst, out_s2828, out_e2828, result2828);
PE P2829(out_s2765, out_e2828, clk, rst, out_s2829, out_e2829, result2829);
PE P2830(out_s2766, out_e2829, clk, rst, out_s2830, out_e2830, result2830);
PE P2831(out_s2767, out_e2830, clk, rst, out_s2831, out_e2831, result2831);
PE P2832(out_s2768, out_e2831, clk, rst, out_s2832, out_e2832, result2832);
PE P2833(out_s2769, out_e2832, clk, rst, out_s2833, out_e2833, result2833);
PE P2834(out_s2770, out_e2833, clk, rst, out_s2834, out_e2834, result2834);
PE P2835(out_s2771, out_e2834, clk, rst, out_s2835, out_e2835, result2835);
PE P2836(out_s2772, out_e2835, clk, rst, out_s2836, out_e2836, result2836);
PE P2837(out_s2773, out_e2836, clk, rst, out_s2837, out_e2837, result2837);
PE P2838(out_s2774, out_e2837, clk, rst, out_s2838, out_e2838, result2838);
PE P2839(out_s2775, out_e2838, clk, rst, out_s2839, out_e2839, result2839);
PE P2840(out_s2776, out_e2839, clk, rst, out_s2840, out_e2840, result2840);
PE P2841(out_s2777, out_e2840, clk, rst, out_s2841, out_e2841, result2841);
PE P2842(out_s2778, out_e2841, clk, rst, out_s2842, out_e2842, result2842);
PE P2843(out_s2779, out_e2842, clk, rst, out_s2843, out_e2843, result2843);
PE P2844(out_s2780, out_e2843, clk, rst, out_s2844, out_e2844, result2844);
PE P2845(out_s2781, out_e2844, clk, rst, out_s2845, out_e2845, result2845);
PE P2846(out_s2782, out_e2845, clk, rst, out_s2846, out_e2846, result2846);
PE P2847(out_s2783, out_e2846, clk, rst, out_s2847, out_e2847, result2847);
PE P2848(out_s2784, out_e2847, clk, rst, out_s2848, out_e2848, result2848);
PE P2849(out_s2785, out_e2848, clk, rst, out_s2849, out_e2849, result2849);
PE P2850(out_s2786, out_e2849, clk, rst, out_s2850, out_e2850, result2850);
PE P2851(out_s2787, out_e2850, clk, rst, out_s2851, out_e2851, result2851);
PE P2852(out_s2788, out_e2851, clk, rst, out_s2852, out_e2852, result2852);
PE P2853(out_s2789, out_e2852, clk, rst, out_s2853, out_e2853, result2853);
PE P2854(out_s2790, out_e2853, clk, rst, out_s2854, out_e2854, result2854);
PE P2855(out_s2791, out_e2854, clk, rst, out_s2855, out_e2855, result2855);
PE P2856(out_s2792, out_e2855, clk, rst, out_s2856, out_e2856, result2856);
PE P2857(out_s2793, out_e2856, clk, rst, out_s2857, out_e2857, result2857);
PE P2858(out_s2794, out_e2857, clk, rst, out_s2858, out_e2858, result2858);
PE P2859(out_s2795, out_e2858, clk, rst, out_s2859, out_e2859, result2859);
PE P2860(out_s2796, out_e2859, clk, rst, out_s2860, out_e2860, result2860);
PE P2861(out_s2797, out_e2860, clk, rst, out_s2861, out_e2861, result2861);
PE P2862(out_s2798, out_e2861, clk, rst, out_s2862, out_e2862, result2862);
PE P2863(out_s2799, out_e2862, clk, rst, out_s2863, out_e2863, result2863);
PE P2864(out_s2800, out_e2863, clk, rst, out_s2864, out_e2864, result2864);
PE P2865(out_s2801, out_e2864, clk, rst, out_s2865, out_e2865, result2865);
PE P2866(out_s2802, out_e2865, clk, rst, out_s2866, out_e2866, result2866);
PE P2867(out_s2803, out_e2866, clk, rst, out_s2867, out_e2867, result2867);
PE P2868(out_s2804, out_e2867, clk, rst, out_s2868, out_e2868, result2868);
PE P2869(out_s2805, out_e2868, clk, rst, out_s2869, out_e2869, result2869);
PE P2870(out_s2806, out_e2869, clk, rst, out_s2870, out_e2870, result2870);
PE P2871(out_s2807, out_e2870, clk, rst, out_s2871, out_e2871, result2871);
PE P2872(out_s2808, out_e2871, clk, rst, out_s2872, out_e2872, result2872);
PE P2873(out_s2809, out_e2872, clk, rst, out_s2873, out_e2873, result2873);
PE P2874(out_s2810, out_e2873, clk, rst, out_s2874, out_e2874, result2874);
PE P2875(out_s2811, out_e2874, clk, rst, out_s2875, out_e2875, result2875);
PE P2876(out_s2812, out_e2875, clk, rst, out_s2876, out_e2876, result2876);
PE P2877(out_s2813, out_e2876, clk, rst, out_s2877, out_e2877, result2877);
PE P2878(out_s2814, out_e2877, clk, rst, out_s2878, out_e2878, result2878);
PE P2879(out_s2815, out_e2878, clk, rst, out_s2879, out_e2879, result2879);

PE P2881(out_s2817, out_e2880, clk, rst, out_s2881, out_e2881, result2881);
PE P2882(out_s2818, out_e2881, clk, rst, out_s2882, out_e2882, result2882);
PE P2883(out_s2819, out_e2882, clk, rst, out_s2883, out_e2883, result2883);
PE P2884(out_s2820, out_e2883, clk, rst, out_s2884, out_e2884, result2884);
PE P2885(out_s2821, out_e2884, clk, rst, out_s2885, out_e2885, result2885);
PE P2886(out_s2822, out_e2885, clk, rst, out_s2886, out_e2886, result2886);
PE P2887(out_s2823, out_e2886, clk, rst, out_s2887, out_e2887, result2887);
PE P2888(out_s2824, out_e2887, clk, rst, out_s2888, out_e2888, result2888);
PE P2889(out_s2825, out_e2888, clk, rst, out_s2889, out_e2889, result2889);
PE P2890(out_s2826, out_e2889, clk, rst, out_s2890, out_e2890, result2890);
PE P2891(out_s2827, out_e2890, clk, rst, out_s2891, out_e2891, result2891);
PE P2892(out_s2828, out_e2891, clk, rst, out_s2892, out_e2892, result2892);
PE P2893(out_s2829, out_e2892, clk, rst, out_s2893, out_e2893, result2893);
PE P2894(out_s2830, out_e2893, clk, rst, out_s2894, out_e2894, result2894);
PE P2895(out_s2831, out_e2894, clk, rst, out_s2895, out_e2895, result2895);
PE P2896(out_s2832, out_e2895, clk, rst, out_s2896, out_e2896, result2896);
PE P2897(out_s2833, out_e2896, clk, rst, out_s2897, out_e2897, result2897);
PE P2898(out_s2834, out_e2897, clk, rst, out_s2898, out_e2898, result2898);
PE P2899(out_s2835, out_e2898, clk, rst, out_s2899, out_e2899, result2899);
PE P2900(out_s2836, out_e2899, clk, rst, out_s2900, out_e2900, result2900);
PE P2901(out_s2837, out_e2900, clk, rst, out_s2901, out_e2901, result2901);
PE P2902(out_s2838, out_e2901, clk, rst, out_s2902, out_e2902, result2902);
PE P2903(out_s2839, out_e2902, clk, rst, out_s2903, out_e2903, result2903);
PE P2904(out_s2840, out_e2903, clk, rst, out_s2904, out_e2904, result2904);
PE P2905(out_s2841, out_e2904, clk, rst, out_s2905, out_e2905, result2905);
PE P2906(out_s2842, out_e2905, clk, rst, out_s2906, out_e2906, result2906);
PE P2907(out_s2843, out_e2906, clk, rst, out_s2907, out_e2907, result2907);
PE P2908(out_s2844, out_e2907, clk, rst, out_s2908, out_e2908, result2908);
PE P2909(out_s2845, out_e2908, clk, rst, out_s2909, out_e2909, result2909);
PE P2910(out_s2846, out_e2909, clk, rst, out_s2910, out_e2910, result2910);
PE P2911(out_s2847, out_e2910, clk, rst, out_s2911, out_e2911, result2911);
PE P2912(out_s2848, out_e2911, clk, rst, out_s2912, out_e2912, result2912);
PE P2913(out_s2849, out_e2912, clk, rst, out_s2913, out_e2913, result2913);
PE P2914(out_s2850, out_e2913, clk, rst, out_s2914, out_e2914, result2914);
PE P2915(out_s2851, out_e2914, clk, rst, out_s2915, out_e2915, result2915);
PE P2916(out_s2852, out_e2915, clk, rst, out_s2916, out_e2916, result2916);
PE P2917(out_s2853, out_e2916, clk, rst, out_s2917, out_e2917, result2917);
PE P2918(out_s2854, out_e2917, clk, rst, out_s2918, out_e2918, result2918);
PE P2919(out_s2855, out_e2918, clk, rst, out_s2919, out_e2919, result2919);
PE P2920(out_s2856, out_e2919, clk, rst, out_s2920, out_e2920, result2920);
PE P2921(out_s2857, out_e2920, clk, rst, out_s2921, out_e2921, result2921);
PE P2922(out_s2858, out_e2921, clk, rst, out_s2922, out_e2922, result2922);
PE P2923(out_s2859, out_e2922, clk, rst, out_s2923, out_e2923, result2923);
PE P2924(out_s2860, out_e2923, clk, rst, out_s2924, out_e2924, result2924);
PE P2925(out_s2861, out_e2924, clk, rst, out_s2925, out_e2925, result2925);
PE P2926(out_s2862, out_e2925, clk, rst, out_s2926, out_e2926, result2926);
PE P2927(out_s2863, out_e2926, clk, rst, out_s2927, out_e2927, result2927);
PE P2928(out_s2864, out_e2927, clk, rst, out_s2928, out_e2928, result2928);
PE P2929(out_s2865, out_e2928, clk, rst, out_s2929, out_e2929, result2929);
PE P2930(out_s2866, out_e2929, clk, rst, out_s2930, out_e2930, result2930);
PE P2931(out_s2867, out_e2930, clk, rst, out_s2931, out_e2931, result2931);
PE P2932(out_s2868, out_e2931, clk, rst, out_s2932, out_e2932, result2932);
PE P2933(out_s2869, out_e2932, clk, rst, out_s2933, out_e2933, result2933);
PE P2934(out_s2870, out_e2933, clk, rst, out_s2934, out_e2934, result2934);
PE P2935(out_s2871, out_e2934, clk, rst, out_s2935, out_e2935, result2935);
PE P2936(out_s2872, out_e2935, clk, rst, out_s2936, out_e2936, result2936);
PE P2937(out_s2873, out_e2936, clk, rst, out_s2937, out_e2937, result2937);
PE P2938(out_s2874, out_e2937, clk, rst, out_s2938, out_e2938, result2938);
PE P2939(out_s2875, out_e2938, clk, rst, out_s2939, out_e2939, result2939);
PE P2940(out_s2876, out_e2939, clk, rst, out_s2940, out_e2940, result2940);
PE P2941(out_s2877, out_e2940, clk, rst, out_s2941, out_e2941, result2941);
PE P2942(out_s2878, out_e2941, clk, rst, out_s2942, out_e2942, result2942);
PE P2943(out_s2879, out_e2942, clk, rst, out_s2943, out_e2943, result2943);

PE P2945(out_s2881, out_e2944, clk, rst, out_s2945, out_e2945, result2945);
PE P2946(out_s2882, out_e2945, clk, rst, out_s2946, out_e2946, result2946);
PE P2947(out_s2883, out_e2946, clk, rst, out_s2947, out_e2947, result2947);
PE P2948(out_s2884, out_e2947, clk, rst, out_s2948, out_e2948, result2948);
PE P2949(out_s2885, out_e2948, clk, rst, out_s2949, out_e2949, result2949);
PE P2950(out_s2886, out_e2949, clk, rst, out_s2950, out_e2950, result2950);
PE P2951(out_s2887, out_e2950, clk, rst, out_s2951, out_e2951, result2951);
PE P2952(out_s2888, out_e2951, clk, rst, out_s2952, out_e2952, result2952);
PE P2953(out_s2889, out_e2952, clk, rst, out_s2953, out_e2953, result2953);
PE P2954(out_s2890, out_e2953, clk, rst, out_s2954, out_e2954, result2954);
PE P2955(out_s2891, out_e2954, clk, rst, out_s2955, out_e2955, result2955);
PE P2956(out_s2892, out_e2955, clk, rst, out_s2956, out_e2956, result2956);
PE P2957(out_s2893, out_e2956, clk, rst, out_s2957, out_e2957, result2957);
PE P2958(out_s2894, out_e2957, clk, rst, out_s2958, out_e2958, result2958);
PE P2959(out_s2895, out_e2958, clk, rst, out_s2959, out_e2959, result2959);
PE P2960(out_s2896, out_e2959, clk, rst, out_s2960, out_e2960, result2960);
PE P2961(out_s2897, out_e2960, clk, rst, out_s2961, out_e2961, result2961);
PE P2962(out_s2898, out_e2961, clk, rst, out_s2962, out_e2962, result2962);
PE P2963(out_s2899, out_e2962, clk, rst, out_s2963, out_e2963, result2963);
PE P2964(out_s2900, out_e2963, clk, rst, out_s2964, out_e2964, result2964);
PE P2965(out_s2901, out_e2964, clk, rst, out_s2965, out_e2965, result2965);
PE P2966(out_s2902, out_e2965, clk, rst, out_s2966, out_e2966, result2966);
PE P2967(out_s2903, out_e2966, clk, rst, out_s2967, out_e2967, result2967);
PE P2968(out_s2904, out_e2967, clk, rst, out_s2968, out_e2968, result2968);
PE P2969(out_s2905, out_e2968, clk, rst, out_s2969, out_e2969, result2969);
PE P2970(out_s2906, out_e2969, clk, rst, out_s2970, out_e2970, result2970);
PE P2971(out_s2907, out_e2970, clk, rst, out_s2971, out_e2971, result2971);
PE P2972(out_s2908, out_e2971, clk, rst, out_s2972, out_e2972, result2972);
PE P2973(out_s2909, out_e2972, clk, rst, out_s2973, out_e2973, result2973);
PE P2974(out_s2910, out_e2973, clk, rst, out_s2974, out_e2974, result2974);
PE P2975(out_s2911, out_e2974, clk, rst, out_s2975, out_e2975, result2975);
PE P2976(out_s2912, out_e2975, clk, rst, out_s2976, out_e2976, result2976);
PE P2977(out_s2913, out_e2976, clk, rst, out_s2977, out_e2977, result2977);
PE P2978(out_s2914, out_e2977, clk, rst, out_s2978, out_e2978, result2978);
PE P2979(out_s2915, out_e2978, clk, rst, out_s2979, out_e2979, result2979);
PE P2980(out_s2916, out_e2979, clk, rst, out_s2980, out_e2980, result2980);
PE P2981(out_s2917, out_e2980, clk, rst, out_s2981, out_e2981, result2981);
PE P2982(out_s2918, out_e2981, clk, rst, out_s2982, out_e2982, result2982);
PE P2983(out_s2919, out_e2982, clk, rst, out_s2983, out_e2983, result2983);
PE P2984(out_s2920, out_e2983, clk, rst, out_s2984, out_e2984, result2984);
PE P2985(out_s2921, out_e2984, clk, rst, out_s2985, out_e2985, result2985);
PE P2986(out_s2922, out_e2985, clk, rst, out_s2986, out_e2986, result2986);
PE P2987(out_s2923, out_e2986, clk, rst, out_s2987, out_e2987, result2987);
PE P2988(out_s2924, out_e2987, clk, rst, out_s2988, out_e2988, result2988);
PE P2989(out_s2925, out_e2988, clk, rst, out_s2989, out_e2989, result2989);
PE P2990(out_s2926, out_e2989, clk, rst, out_s2990, out_e2990, result2990);
PE P2991(out_s2927, out_e2990, clk, rst, out_s2991, out_e2991, result2991);
PE P2992(out_s2928, out_e2991, clk, rst, out_s2992, out_e2992, result2992);
PE P2993(out_s2929, out_e2992, clk, rst, out_s2993, out_e2993, result2993);
PE P2994(out_s2930, out_e2993, clk, rst, out_s2994, out_e2994, result2994);
PE P2995(out_s2931, out_e2994, clk, rst, out_s2995, out_e2995, result2995);
PE P2996(out_s2932, out_e2995, clk, rst, out_s2996, out_e2996, result2996);
PE P2997(out_s2933, out_e2996, clk, rst, out_s2997, out_e2997, result2997);
PE P2998(out_s2934, out_e2997, clk, rst, out_s2998, out_e2998, result2998);
PE P2999(out_s2935, out_e2998, clk, rst, out_s2999, out_e2999, result2999);
PE P3000(out_s2936, out_e2999, clk, rst, out_s3000, out_e3000, result3000);
PE P3001(out_s2937, out_e3000, clk, rst, out_s3001, out_e3001, result3001);
PE P3002(out_s2938, out_e3001, clk, rst, out_s3002, out_e3002, result3002);
PE P3003(out_s2939, out_e3002, clk, rst, out_s3003, out_e3003, result3003);
PE P3004(out_s2940, out_e3003, clk, rst, out_s3004, out_e3004, result3004);
PE P3005(out_s2941, out_e3004, clk, rst, out_s3005, out_e3005, result3005);
PE P3006(out_s2942, out_e3005, clk, rst, out_s3006, out_e3006, result3006);
PE P3007(out_s2943, out_e3006, clk, rst, out_s3007, out_e3007, result3007);

PE P3009(out_s2945, out_e3008, clk, rst, out_s3009, out_e3009, result3009);
PE P3010(out_s2946, out_e3009, clk, rst, out_s3010, out_e3010, result3010);
PE P3011(out_s2947, out_e3010, clk, rst, out_s3011, out_e3011, result3011);
PE P3012(out_s2948, out_e3011, clk, rst, out_s3012, out_e3012, result3012);
PE P3013(out_s2949, out_e3012, clk, rst, out_s3013, out_e3013, result3013);
PE P3014(out_s2950, out_e3013, clk, rst, out_s3014, out_e3014, result3014);
PE P3015(out_s2951, out_e3014, clk, rst, out_s3015, out_e3015, result3015);
PE P3016(out_s2952, out_e3015, clk, rst, out_s3016, out_e3016, result3016);
PE P3017(out_s2953, out_e3016, clk, rst, out_s3017, out_e3017, result3017);
PE P3018(out_s2954, out_e3017, clk, rst, out_s3018, out_e3018, result3018);
PE P3019(out_s2955, out_e3018, clk, rst, out_s3019, out_e3019, result3019);
PE P3020(out_s2956, out_e3019, clk, rst, out_s3020, out_e3020, result3020);
PE P3021(out_s2957, out_e3020, clk, rst, out_s3021, out_e3021, result3021);
PE P3022(out_s2958, out_e3021, clk, rst, out_s3022, out_e3022, result3022);
PE P3023(out_s2959, out_e3022, clk, rst, out_s3023, out_e3023, result3023);
PE P3024(out_s2960, out_e3023, clk, rst, out_s3024, out_e3024, result3024);
PE P3025(out_s2961, out_e3024, clk, rst, out_s3025, out_e3025, result3025);
PE P3026(out_s2962, out_e3025, clk, rst, out_s3026, out_e3026, result3026);
PE P3027(out_s2963, out_e3026, clk, rst, out_s3027, out_e3027, result3027);
PE P3028(out_s2964, out_e3027, clk, rst, out_s3028, out_e3028, result3028);
PE P3029(out_s2965, out_e3028, clk, rst, out_s3029, out_e3029, result3029);
PE P3030(out_s2966, out_e3029, clk, rst, out_s3030, out_e3030, result3030);
PE P3031(out_s2967, out_e3030, clk, rst, out_s3031, out_e3031, result3031);
PE P3032(out_s2968, out_e3031, clk, rst, out_s3032, out_e3032, result3032);
PE P3033(out_s2969, out_e3032, clk, rst, out_s3033, out_e3033, result3033);
PE P3034(out_s2970, out_e3033, clk, rst, out_s3034, out_e3034, result3034);
PE P3035(out_s2971, out_e3034, clk, rst, out_s3035, out_e3035, result3035);
PE P3036(out_s2972, out_e3035, clk, rst, out_s3036, out_e3036, result3036);
PE P3037(out_s2973, out_e3036, clk, rst, out_s3037, out_e3037, result3037);
PE P3038(out_s2974, out_e3037, clk, rst, out_s3038, out_e3038, result3038);
PE P3039(out_s2975, out_e3038, clk, rst, out_s3039, out_e3039, result3039);
PE P3040(out_s2976, out_e3039, clk, rst, out_s3040, out_e3040, result3040);
PE P3041(out_s2977, out_e3040, clk, rst, out_s3041, out_e3041, result3041);
PE P3042(out_s2978, out_e3041, clk, rst, out_s3042, out_e3042, result3042);
PE P3043(out_s2979, out_e3042, clk, rst, out_s3043, out_e3043, result3043);
PE P3044(out_s2980, out_e3043, clk, rst, out_s3044, out_e3044, result3044);
PE P3045(out_s2981, out_e3044, clk, rst, out_s3045, out_e3045, result3045);
PE P3046(out_s2982, out_e3045, clk, rst, out_s3046, out_e3046, result3046);
PE P3047(out_s2983, out_e3046, clk, rst, out_s3047, out_e3047, result3047);
PE P3048(out_s2984, out_e3047, clk, rst, out_s3048, out_e3048, result3048);
PE P3049(out_s2985, out_e3048, clk, rst, out_s3049, out_e3049, result3049);
PE P3050(out_s2986, out_e3049, clk, rst, out_s3050, out_e3050, result3050);
PE P3051(out_s2987, out_e3050, clk, rst, out_s3051, out_e3051, result3051);
PE P3052(out_s2988, out_e3051, clk, rst, out_s3052, out_e3052, result3052);
PE P3053(out_s2989, out_e3052, clk, rst, out_s3053, out_e3053, result3053);
PE P3054(out_s2990, out_e3053, clk, rst, out_s3054, out_e3054, result3054);
PE P3055(out_s2991, out_e3054, clk, rst, out_s3055, out_e3055, result3055);
PE P3056(out_s2992, out_e3055, clk, rst, out_s3056, out_e3056, result3056);
PE P3057(out_s2993, out_e3056, clk, rst, out_s3057, out_e3057, result3057);
PE P3058(out_s2994, out_e3057, clk, rst, out_s3058, out_e3058, result3058);
PE P3059(out_s2995, out_e3058, clk, rst, out_s3059, out_e3059, result3059);
PE P3060(out_s2996, out_e3059, clk, rst, out_s3060, out_e3060, result3060);
PE P3061(out_s2997, out_e3060, clk, rst, out_s3061, out_e3061, result3061);
PE P3062(out_s2998, out_e3061, clk, rst, out_s3062, out_e3062, result3062);
PE P3063(out_s2999, out_e3062, clk, rst, out_s3063, out_e3063, result3063);
PE P3064(out_s3000, out_e3063, clk, rst, out_s3064, out_e3064, result3064);
PE P3065(out_s3001, out_e3064, clk, rst, out_s3065, out_e3065, result3065);
PE P3066(out_s3002, out_e3065, clk, rst, out_s3066, out_e3066, result3066);
PE P3067(out_s3003, out_e3066, clk, rst, out_s3067, out_e3067, result3067);
PE P3068(out_s3004, out_e3067, clk, rst, out_s3068, out_e3068, result3068);
PE P3069(out_s3005, out_e3068, clk, rst, out_s3069, out_e3069, result3069);
PE P3070(out_s3006, out_e3069, clk, rst, out_s3070, out_e3070, result3070);
PE P3071(out_s3007, out_e3070, clk, rst, out_s3071, out_e3071, result3071);

PE P3073(out_s3009, out_e3072, clk, rst, out_s3073, out_e3073, result3073);
PE P3074(out_s3010, out_e3073, clk, rst, out_s3074, out_e3074, result3074);
PE P3075(out_s3011, out_e3074, clk, rst, out_s3075, out_e3075, result3075);
PE P3076(out_s3012, out_e3075, clk, rst, out_s3076, out_e3076, result3076);
PE P3077(out_s3013, out_e3076, clk, rst, out_s3077, out_e3077, result3077);
PE P3078(out_s3014, out_e3077, clk, rst, out_s3078, out_e3078, result3078);
PE P3079(out_s3015, out_e3078, clk, rst, out_s3079, out_e3079, result3079);
PE P3080(out_s3016, out_e3079, clk, rst, out_s3080, out_e3080, result3080);
PE P3081(out_s3017, out_e3080, clk, rst, out_s3081, out_e3081, result3081);
PE P3082(out_s3018, out_e3081, clk, rst, out_s3082, out_e3082, result3082);
PE P3083(out_s3019, out_e3082, clk, rst, out_s3083, out_e3083, result3083);
PE P3084(out_s3020, out_e3083, clk, rst, out_s3084, out_e3084, result3084);
PE P3085(out_s3021, out_e3084, clk, rst, out_s3085, out_e3085, result3085);
PE P3086(out_s3022, out_e3085, clk, rst, out_s3086, out_e3086, result3086);
PE P3087(out_s3023, out_e3086, clk, rst, out_s3087, out_e3087, result3087);
PE P3088(out_s3024, out_e3087, clk, rst, out_s3088, out_e3088, result3088);
PE P3089(out_s3025, out_e3088, clk, rst, out_s3089, out_e3089, result3089);
PE P3090(out_s3026, out_e3089, clk, rst, out_s3090, out_e3090, result3090);
PE P3091(out_s3027, out_e3090, clk, rst, out_s3091, out_e3091, result3091);
PE P3092(out_s3028, out_e3091, clk, rst, out_s3092, out_e3092, result3092);
PE P3093(out_s3029, out_e3092, clk, rst, out_s3093, out_e3093, result3093);
PE P3094(out_s3030, out_e3093, clk, rst, out_s3094, out_e3094, result3094);
PE P3095(out_s3031, out_e3094, clk, rst, out_s3095, out_e3095, result3095);
PE P3096(out_s3032, out_e3095, clk, rst, out_s3096, out_e3096, result3096);
PE P3097(out_s3033, out_e3096, clk, rst, out_s3097, out_e3097, result3097);
PE P3098(out_s3034, out_e3097, clk, rst, out_s3098, out_e3098, result3098);
PE P3099(out_s3035, out_e3098, clk, rst, out_s3099, out_e3099, result3099);
PE P3100(out_s3036, out_e3099, clk, rst, out_s3100, out_e3100, result3100);
PE P3101(out_s3037, out_e3100, clk, rst, out_s3101, out_e3101, result3101);
PE P3102(out_s3038, out_e3101, clk, rst, out_s3102, out_e3102, result3102);
PE P3103(out_s3039, out_e3102, clk, rst, out_s3103, out_e3103, result3103);
PE P3104(out_s3040, out_e3103, clk, rst, out_s3104, out_e3104, result3104);
PE P3105(out_s3041, out_e3104, clk, rst, out_s3105, out_e3105, result3105);
PE P3106(out_s3042, out_e3105, clk, rst, out_s3106, out_e3106, result3106);
PE P3107(out_s3043, out_e3106, clk, rst, out_s3107, out_e3107, result3107);
PE P3108(out_s3044, out_e3107, clk, rst, out_s3108, out_e3108, result3108);
PE P3109(out_s3045, out_e3108, clk, rst, out_s3109, out_e3109, result3109);
PE P3110(out_s3046, out_e3109, clk, rst, out_s3110, out_e3110, result3110);
PE P3111(out_s3047, out_e3110, clk, rst, out_s3111, out_e3111, result3111);
PE P3112(out_s3048, out_e3111, clk, rst, out_s3112, out_e3112, result3112);
PE P3113(out_s3049, out_e3112, clk, rst, out_s3113, out_e3113, result3113);
PE P3114(out_s3050, out_e3113, clk, rst, out_s3114, out_e3114, result3114);
PE P3115(out_s3051, out_e3114, clk, rst, out_s3115, out_e3115, result3115);
PE P3116(out_s3052, out_e3115, clk, rst, out_s3116, out_e3116, result3116);
PE P3117(out_s3053, out_e3116, clk, rst, out_s3117, out_e3117, result3117);
PE P3118(out_s3054, out_e3117, clk, rst, out_s3118, out_e3118, result3118);
PE P3119(out_s3055, out_e3118, clk, rst, out_s3119, out_e3119, result3119);
PE P3120(out_s3056, out_e3119, clk, rst, out_s3120, out_e3120, result3120);
PE P3121(out_s3057, out_e3120, clk, rst, out_s3121, out_e3121, result3121);
PE P3122(out_s3058, out_e3121, clk, rst, out_s3122, out_e3122, result3122);
PE P3123(out_s3059, out_e3122, clk, rst, out_s3123, out_e3123, result3123);
PE P3124(out_s3060, out_e3123, clk, rst, out_s3124, out_e3124, result3124);
PE P3125(out_s3061, out_e3124, clk, rst, out_s3125, out_e3125, result3125);
PE P3126(out_s3062, out_e3125, clk, rst, out_s3126, out_e3126, result3126);
PE P3127(out_s3063, out_e3126, clk, rst, out_s3127, out_e3127, result3127);
PE P3128(out_s3064, out_e3127, clk, rst, out_s3128, out_e3128, result3128);
PE P3129(out_s3065, out_e3128, clk, rst, out_s3129, out_e3129, result3129);
PE P3130(out_s3066, out_e3129, clk, rst, out_s3130, out_e3130, result3130);
PE P3131(out_s3067, out_e3130, clk, rst, out_s3131, out_e3131, result3131);
PE P3132(out_s3068, out_e3131, clk, rst, out_s3132, out_e3132, result3132);
PE P3133(out_s3069, out_e3132, clk, rst, out_s3133, out_e3133, result3133);
PE P3134(out_s3070, out_e3133, clk, rst, out_s3134, out_e3134, result3134);
PE P3135(out_s3071, out_e3134, clk, rst, out_s3135, out_e3135, result3135);

PE P3137(out_s3073, out_e3136, clk, rst, out_s3137, out_e3137, result3137);
PE P3138(out_s3074, out_e3137, clk, rst, out_s3138, out_e3138, result3138);
PE P3139(out_s3075, out_e3138, clk, rst, out_s3139, out_e3139, result3139);
PE P3140(out_s3076, out_e3139, clk, rst, out_s3140, out_e3140, result3140);
PE P3141(out_s3077, out_e3140, clk, rst, out_s3141, out_e3141, result3141);
PE P3142(out_s3078, out_e3141, clk, rst, out_s3142, out_e3142, result3142);
PE P3143(out_s3079, out_e3142, clk, rst, out_s3143, out_e3143, result3143);
PE P3144(out_s3080, out_e3143, clk, rst, out_s3144, out_e3144, result3144);
PE P3145(out_s3081, out_e3144, clk, rst, out_s3145, out_e3145, result3145);
PE P3146(out_s3082, out_e3145, clk, rst, out_s3146, out_e3146, result3146);
PE P3147(out_s3083, out_e3146, clk, rst, out_s3147, out_e3147, result3147);
PE P3148(out_s3084, out_e3147, clk, rst, out_s3148, out_e3148, result3148);
PE P3149(out_s3085, out_e3148, clk, rst, out_s3149, out_e3149, result3149);
PE P3150(out_s3086, out_e3149, clk, rst, out_s3150, out_e3150, result3150);
PE P3151(out_s3087, out_e3150, clk, rst, out_s3151, out_e3151, result3151);
PE P3152(out_s3088, out_e3151, clk, rst, out_s3152, out_e3152, result3152);
PE P3153(out_s3089, out_e3152, clk, rst, out_s3153, out_e3153, result3153);
PE P3154(out_s3090, out_e3153, clk, rst, out_s3154, out_e3154, result3154);
PE P3155(out_s3091, out_e3154, clk, rst, out_s3155, out_e3155, result3155);
PE P3156(out_s3092, out_e3155, clk, rst, out_s3156, out_e3156, result3156);
PE P3157(out_s3093, out_e3156, clk, rst, out_s3157, out_e3157, result3157);
PE P3158(out_s3094, out_e3157, clk, rst, out_s3158, out_e3158, result3158);
PE P3159(out_s3095, out_e3158, clk, rst, out_s3159, out_e3159, result3159);
PE P3160(out_s3096, out_e3159, clk, rst, out_s3160, out_e3160, result3160);
PE P3161(out_s3097, out_e3160, clk, rst, out_s3161, out_e3161, result3161);
PE P3162(out_s3098, out_e3161, clk, rst, out_s3162, out_e3162, result3162);
PE P3163(out_s3099, out_e3162, clk, rst, out_s3163, out_e3163, result3163);
PE P3164(out_s3100, out_e3163, clk, rst, out_s3164, out_e3164, result3164);
PE P3165(out_s3101, out_e3164, clk, rst, out_s3165, out_e3165, result3165);
PE P3166(out_s3102, out_e3165, clk, rst, out_s3166, out_e3166, result3166);
PE P3167(out_s3103, out_e3166, clk, rst, out_s3167, out_e3167, result3167);
PE P3168(out_s3104, out_e3167, clk, rst, out_s3168, out_e3168, result3168);
PE P3169(out_s3105, out_e3168, clk, rst, out_s3169, out_e3169, result3169);
PE P3170(out_s3106, out_e3169, clk, rst, out_s3170, out_e3170, result3170);
PE P3171(out_s3107, out_e3170, clk, rst, out_s3171, out_e3171, result3171);
PE P3172(out_s3108, out_e3171, clk, rst, out_s3172, out_e3172, result3172);
PE P3173(out_s3109, out_e3172, clk, rst, out_s3173, out_e3173, result3173);
PE P3174(out_s3110, out_e3173, clk, rst, out_s3174, out_e3174, result3174);
PE P3175(out_s3111, out_e3174, clk, rst, out_s3175, out_e3175, result3175);
PE P3176(out_s3112, out_e3175, clk, rst, out_s3176, out_e3176, result3176);
PE P3177(out_s3113, out_e3176, clk, rst, out_s3177, out_e3177, result3177);
PE P3178(out_s3114, out_e3177, clk, rst, out_s3178, out_e3178, result3178);
PE P3179(out_s3115, out_e3178, clk, rst, out_s3179, out_e3179, result3179);
PE P3180(out_s3116, out_e3179, clk, rst, out_s3180, out_e3180, result3180);
PE P3181(out_s3117, out_e3180, clk, rst, out_s3181, out_e3181, result3181);
PE P3182(out_s3118, out_e3181, clk, rst, out_s3182, out_e3182, result3182);
PE P3183(out_s3119, out_e3182, clk, rst, out_s3183, out_e3183, result3183);
PE P3184(out_s3120, out_e3183, clk, rst, out_s3184, out_e3184, result3184);
PE P3185(out_s3121, out_e3184, clk, rst, out_s3185, out_e3185, result3185);
PE P3186(out_s3122, out_e3185, clk, rst, out_s3186, out_e3186, result3186);
PE P3187(out_s3123, out_e3186, clk, rst, out_s3187, out_e3187, result3187);
PE P3188(out_s3124, out_e3187, clk, rst, out_s3188, out_e3188, result3188);
PE P3189(out_s3125, out_e3188, clk, rst, out_s3189, out_e3189, result3189);
PE P3190(out_s3126, out_e3189, clk, rst, out_s3190, out_e3190, result3190);
PE P3191(out_s3127, out_e3190, clk, rst, out_s3191, out_e3191, result3191);
PE P3192(out_s3128, out_e3191, clk, rst, out_s3192, out_e3192, result3192);
PE P3193(out_s3129, out_e3192, clk, rst, out_s3193, out_e3193, result3193);
PE P3194(out_s3130, out_e3193, clk, rst, out_s3194, out_e3194, result3194);
PE P3195(out_s3131, out_e3194, clk, rst, out_s3195, out_e3195, result3195);
PE P3196(out_s3132, out_e3195, clk, rst, out_s3196, out_e3196, result3196);
PE P3197(out_s3133, out_e3196, clk, rst, out_s3197, out_e3197, result3197);
PE P3198(out_s3134, out_e3197, clk, rst, out_s3198, out_e3198, result3198);
PE P3199(out_s3135, out_e3198, clk, rst, out_s3199, out_e3199, result3199);

PE P3201(out_s3137, out_e3200, clk, rst, out_s3201, out_e3201, result3201);
PE P3202(out_s3138, out_e3201, clk, rst, out_s3202, out_e3202, result3202);
PE P3203(out_s3139, out_e3202, clk, rst, out_s3203, out_e3203, result3203);
PE P3204(out_s3140, out_e3203, clk, rst, out_s3204, out_e3204, result3204);
PE P3205(out_s3141, out_e3204, clk, rst, out_s3205, out_e3205, result3205);
PE P3206(out_s3142, out_e3205, clk, rst, out_s3206, out_e3206, result3206);
PE P3207(out_s3143, out_e3206, clk, rst, out_s3207, out_e3207, result3207);
PE P3208(out_s3144, out_e3207, clk, rst, out_s3208, out_e3208, result3208);
PE P3209(out_s3145, out_e3208, clk, rst, out_s3209, out_e3209, result3209);
PE P3210(out_s3146, out_e3209, clk, rst, out_s3210, out_e3210, result3210);
PE P3211(out_s3147, out_e3210, clk, rst, out_s3211, out_e3211, result3211);
PE P3212(out_s3148, out_e3211, clk, rst, out_s3212, out_e3212, result3212);
PE P3213(out_s3149, out_e3212, clk, rst, out_s3213, out_e3213, result3213);
PE P3214(out_s3150, out_e3213, clk, rst, out_s3214, out_e3214, result3214);
PE P3215(out_s3151, out_e3214, clk, rst, out_s3215, out_e3215, result3215);
PE P3216(out_s3152, out_e3215, clk, rst, out_s3216, out_e3216, result3216);
PE P3217(out_s3153, out_e3216, clk, rst, out_s3217, out_e3217, result3217);
PE P3218(out_s3154, out_e3217, clk, rst, out_s3218, out_e3218, result3218);
PE P3219(out_s3155, out_e3218, clk, rst, out_s3219, out_e3219, result3219);
PE P3220(out_s3156, out_e3219, clk, rst, out_s3220, out_e3220, result3220);
PE P3221(out_s3157, out_e3220, clk, rst, out_s3221, out_e3221, result3221);
PE P3222(out_s3158, out_e3221, clk, rst, out_s3222, out_e3222, result3222);
PE P3223(out_s3159, out_e3222, clk, rst, out_s3223, out_e3223, result3223);
PE P3224(out_s3160, out_e3223, clk, rst, out_s3224, out_e3224, result3224);
PE P3225(out_s3161, out_e3224, clk, rst, out_s3225, out_e3225, result3225);
PE P3226(out_s3162, out_e3225, clk, rst, out_s3226, out_e3226, result3226);
PE P3227(out_s3163, out_e3226, clk, rst, out_s3227, out_e3227, result3227);
PE P3228(out_s3164, out_e3227, clk, rst, out_s3228, out_e3228, result3228);
PE P3229(out_s3165, out_e3228, clk, rst, out_s3229, out_e3229, result3229);
PE P3230(out_s3166, out_e3229, clk, rst, out_s3230, out_e3230, result3230);
PE P3231(out_s3167, out_e3230, clk, rst, out_s3231, out_e3231, result3231);
PE P3232(out_s3168, out_e3231, clk, rst, out_s3232, out_e3232, result3232);
PE P3233(out_s3169, out_e3232, clk, rst, out_s3233, out_e3233, result3233);
PE P3234(out_s3170, out_e3233, clk, rst, out_s3234, out_e3234, result3234);
PE P3235(out_s3171, out_e3234, clk, rst, out_s3235, out_e3235, result3235);
PE P3236(out_s3172, out_e3235, clk, rst, out_s3236, out_e3236, result3236);
PE P3237(out_s3173, out_e3236, clk, rst, out_s3237, out_e3237, result3237);
PE P3238(out_s3174, out_e3237, clk, rst, out_s3238, out_e3238, result3238);
PE P3239(out_s3175, out_e3238, clk, rst, out_s3239, out_e3239, result3239);
PE P3240(out_s3176, out_e3239, clk, rst, out_s3240, out_e3240, result3240);
PE P3241(out_s3177, out_e3240, clk, rst, out_s3241, out_e3241, result3241);
PE P3242(out_s3178, out_e3241, clk, rst, out_s3242, out_e3242, result3242);
PE P3243(out_s3179, out_e3242, clk, rst, out_s3243, out_e3243, result3243);
PE P3244(out_s3180, out_e3243, clk, rst, out_s3244, out_e3244, result3244);
PE P3245(out_s3181, out_e3244, clk, rst, out_s3245, out_e3245, result3245);
PE P3246(out_s3182, out_e3245, clk, rst, out_s3246, out_e3246, result3246);
PE P3247(out_s3183, out_e3246, clk, rst, out_s3247, out_e3247, result3247);
PE P3248(out_s3184, out_e3247, clk, rst, out_s3248, out_e3248, result3248);
PE P3249(out_s3185, out_e3248, clk, rst, out_s3249, out_e3249, result3249);
PE P3250(out_s3186, out_e3249, clk, rst, out_s3250, out_e3250, result3250);
PE P3251(out_s3187, out_e3250, clk, rst, out_s3251, out_e3251, result3251);
PE P3252(out_s3188, out_e3251, clk, rst, out_s3252, out_e3252, result3252);
PE P3253(out_s3189, out_e3252, clk, rst, out_s3253, out_e3253, result3253);
PE P3254(out_s3190, out_e3253, clk, rst, out_s3254, out_e3254, result3254);
PE P3255(out_s3191, out_e3254, clk, rst, out_s3255, out_e3255, result3255);
PE P3256(out_s3192, out_e3255, clk, rst, out_s3256, out_e3256, result3256);
PE P3257(out_s3193, out_e3256, clk, rst, out_s3257, out_e3257, result3257);
PE P3258(out_s3194, out_e3257, clk, rst, out_s3258, out_e3258, result3258);
PE P3259(out_s3195, out_e3258, clk, rst, out_s3259, out_e3259, result3259);
PE P3260(out_s3196, out_e3259, clk, rst, out_s3260, out_e3260, result3260);
PE P3261(out_s3197, out_e3260, clk, rst, out_s3261, out_e3261, result3261);
PE P3262(out_s3198, out_e3261, clk, rst, out_s3262, out_e3262, result3262);
PE P3263(out_s3199, out_e3262, clk, rst, out_s3263, out_e3263, result3263);

PE P3265(out_s3201, out_e3264, clk, rst, out_s3265, out_e3265, result3265);
PE P3266(out_s3202, out_e3265, clk, rst, out_s3266, out_e3266, result3266);
PE P3267(out_s3203, out_e3266, clk, rst, out_s3267, out_e3267, result3267);
PE P3268(out_s3204, out_e3267, clk, rst, out_s3268, out_e3268, result3268);
PE P3269(out_s3205, out_e3268, clk, rst, out_s3269, out_e3269, result3269);
PE P3270(out_s3206, out_e3269, clk, rst, out_s3270, out_e3270, result3270);
PE P3271(out_s3207, out_e3270, clk, rst, out_s3271, out_e3271, result3271);
PE P3272(out_s3208, out_e3271, clk, rst, out_s3272, out_e3272, result3272);
PE P3273(out_s3209, out_e3272, clk, rst, out_s3273, out_e3273, result3273);
PE P3274(out_s3210, out_e3273, clk, rst, out_s3274, out_e3274, result3274);
PE P3275(out_s3211, out_e3274, clk, rst, out_s3275, out_e3275, result3275);
PE P3276(out_s3212, out_e3275, clk, rst, out_s3276, out_e3276, result3276);
PE P3277(out_s3213, out_e3276, clk, rst, out_s3277, out_e3277, result3277);
PE P3278(out_s3214, out_e3277, clk, rst, out_s3278, out_e3278, result3278);
PE P3279(out_s3215, out_e3278, clk, rst, out_s3279, out_e3279, result3279);
PE P3280(out_s3216, out_e3279, clk, rst, out_s3280, out_e3280, result3280);
PE P3281(out_s3217, out_e3280, clk, rst, out_s3281, out_e3281, result3281);
PE P3282(out_s3218, out_e3281, clk, rst, out_s3282, out_e3282, result3282);
PE P3283(out_s3219, out_e3282, clk, rst, out_s3283, out_e3283, result3283);
PE P3284(out_s3220, out_e3283, clk, rst, out_s3284, out_e3284, result3284);
PE P3285(out_s3221, out_e3284, clk, rst, out_s3285, out_e3285, result3285);
PE P3286(out_s3222, out_e3285, clk, rst, out_s3286, out_e3286, result3286);
PE P3287(out_s3223, out_e3286, clk, rst, out_s3287, out_e3287, result3287);
PE P3288(out_s3224, out_e3287, clk, rst, out_s3288, out_e3288, result3288);
PE P3289(out_s3225, out_e3288, clk, rst, out_s3289, out_e3289, result3289);
PE P3290(out_s3226, out_e3289, clk, rst, out_s3290, out_e3290, result3290);
PE P3291(out_s3227, out_e3290, clk, rst, out_s3291, out_e3291, result3291);
PE P3292(out_s3228, out_e3291, clk, rst, out_s3292, out_e3292, result3292);
PE P3293(out_s3229, out_e3292, clk, rst, out_s3293, out_e3293, result3293);
PE P3294(out_s3230, out_e3293, clk, rst, out_s3294, out_e3294, result3294);
PE P3295(out_s3231, out_e3294, clk, rst, out_s3295, out_e3295, result3295);
PE P3296(out_s3232, out_e3295, clk, rst, out_s3296, out_e3296, result3296);
PE P3297(out_s3233, out_e3296, clk, rst, out_s3297, out_e3297, result3297);
PE P3298(out_s3234, out_e3297, clk, rst, out_s3298, out_e3298, result3298);
PE P3299(out_s3235, out_e3298, clk, rst, out_s3299, out_e3299, result3299);
PE P3300(out_s3236, out_e3299, clk, rst, out_s3300, out_e3300, result3300);
PE P3301(out_s3237, out_e3300, clk, rst, out_s3301, out_e3301, result3301);
PE P3302(out_s3238, out_e3301, clk, rst, out_s3302, out_e3302, result3302);
PE P3303(out_s3239, out_e3302, clk, rst, out_s3303, out_e3303, result3303);
PE P3304(out_s3240, out_e3303, clk, rst, out_s3304, out_e3304, result3304);
PE P3305(out_s3241, out_e3304, clk, rst, out_s3305, out_e3305, result3305);
PE P3306(out_s3242, out_e3305, clk, rst, out_s3306, out_e3306, result3306);
PE P3307(out_s3243, out_e3306, clk, rst, out_s3307, out_e3307, result3307);
PE P3308(out_s3244, out_e3307, clk, rst, out_s3308, out_e3308, result3308);
PE P3309(out_s3245, out_e3308, clk, rst, out_s3309, out_e3309, result3309);
PE P3310(out_s3246, out_e3309, clk, rst, out_s3310, out_e3310, result3310);
PE P3311(out_s3247, out_e3310, clk, rst, out_s3311, out_e3311, result3311);
PE P3312(out_s3248, out_e3311, clk, rst, out_s3312, out_e3312, result3312);
PE P3313(out_s3249, out_e3312, clk, rst, out_s3313, out_e3313, result3313);
PE P3314(out_s3250, out_e3313, clk, rst, out_s3314, out_e3314, result3314);
PE P3315(out_s3251, out_e3314, clk, rst, out_s3315, out_e3315, result3315);
PE P3316(out_s3252, out_e3315, clk, rst, out_s3316, out_e3316, result3316);
PE P3317(out_s3253, out_e3316, clk, rst, out_s3317, out_e3317, result3317);
PE P3318(out_s3254, out_e3317, clk, rst, out_s3318, out_e3318, result3318);
PE P3319(out_s3255, out_e3318, clk, rst, out_s3319, out_e3319, result3319);
PE P3320(out_s3256, out_e3319, clk, rst, out_s3320, out_e3320, result3320);
PE P3321(out_s3257, out_e3320, clk, rst, out_s3321, out_e3321, result3321);
PE P3322(out_s3258, out_e3321, clk, rst, out_s3322, out_e3322, result3322);
PE P3323(out_s3259, out_e3322, clk, rst, out_s3323, out_e3323, result3323);
PE P3324(out_s3260, out_e3323, clk, rst, out_s3324, out_e3324, result3324);
PE P3325(out_s3261, out_e3324, clk, rst, out_s3325, out_e3325, result3325);
PE P3326(out_s3262, out_e3325, clk, rst, out_s3326, out_e3326, result3326);
PE P3327(out_s3263, out_e3326, clk, rst, out_s3327, out_e3327, result3327);

PE P3329(out_s3265, out_e3328, clk, rst, out_s3329, out_e3329, result3329);
PE P3330(out_s3266, out_e3329, clk, rst, out_s3330, out_e3330, result3330);
PE P3331(out_s3267, out_e3330, clk, rst, out_s3331, out_e3331, result3331);
PE P3332(out_s3268, out_e3331, clk, rst, out_s3332, out_e3332, result3332);
PE P3333(out_s3269, out_e3332, clk, rst, out_s3333, out_e3333, result3333);
PE P3334(out_s3270, out_e3333, clk, rst, out_s3334, out_e3334, result3334);
PE P3335(out_s3271, out_e3334, clk, rst, out_s3335, out_e3335, result3335);
PE P3336(out_s3272, out_e3335, clk, rst, out_s3336, out_e3336, result3336);
PE P3337(out_s3273, out_e3336, clk, rst, out_s3337, out_e3337, result3337);
PE P3338(out_s3274, out_e3337, clk, rst, out_s3338, out_e3338, result3338);
PE P3339(out_s3275, out_e3338, clk, rst, out_s3339, out_e3339, result3339);
PE P3340(out_s3276, out_e3339, clk, rst, out_s3340, out_e3340, result3340);
PE P3341(out_s3277, out_e3340, clk, rst, out_s3341, out_e3341, result3341);
PE P3342(out_s3278, out_e3341, clk, rst, out_s3342, out_e3342, result3342);
PE P3343(out_s3279, out_e3342, clk, rst, out_s3343, out_e3343, result3343);
PE P3344(out_s3280, out_e3343, clk, rst, out_s3344, out_e3344, result3344);
PE P3345(out_s3281, out_e3344, clk, rst, out_s3345, out_e3345, result3345);
PE P3346(out_s3282, out_e3345, clk, rst, out_s3346, out_e3346, result3346);
PE P3347(out_s3283, out_e3346, clk, rst, out_s3347, out_e3347, result3347);
PE P3348(out_s3284, out_e3347, clk, rst, out_s3348, out_e3348, result3348);
PE P3349(out_s3285, out_e3348, clk, rst, out_s3349, out_e3349, result3349);
PE P3350(out_s3286, out_e3349, clk, rst, out_s3350, out_e3350, result3350);
PE P3351(out_s3287, out_e3350, clk, rst, out_s3351, out_e3351, result3351);
PE P3352(out_s3288, out_e3351, clk, rst, out_s3352, out_e3352, result3352);
PE P3353(out_s3289, out_e3352, clk, rst, out_s3353, out_e3353, result3353);
PE P3354(out_s3290, out_e3353, clk, rst, out_s3354, out_e3354, result3354);
PE P3355(out_s3291, out_e3354, clk, rst, out_s3355, out_e3355, result3355);
PE P3356(out_s3292, out_e3355, clk, rst, out_s3356, out_e3356, result3356);
PE P3357(out_s3293, out_e3356, clk, rst, out_s3357, out_e3357, result3357);
PE P3358(out_s3294, out_e3357, clk, rst, out_s3358, out_e3358, result3358);
PE P3359(out_s3295, out_e3358, clk, rst, out_s3359, out_e3359, result3359);
PE P3360(out_s3296, out_e3359, clk, rst, out_s3360, out_e3360, result3360);
PE P3361(out_s3297, out_e3360, clk, rst, out_s3361, out_e3361, result3361);
PE P3362(out_s3298, out_e3361, clk, rst, out_s3362, out_e3362, result3362);
PE P3363(out_s3299, out_e3362, clk, rst, out_s3363, out_e3363, result3363);
PE P3364(out_s3300, out_e3363, clk, rst, out_s3364, out_e3364, result3364);
PE P3365(out_s3301, out_e3364, clk, rst, out_s3365, out_e3365, result3365);
PE P3366(out_s3302, out_e3365, clk, rst, out_s3366, out_e3366, result3366);
PE P3367(out_s3303, out_e3366, clk, rst, out_s3367, out_e3367, result3367);
PE P3368(out_s3304, out_e3367, clk, rst, out_s3368, out_e3368, result3368);
PE P3369(out_s3305, out_e3368, clk, rst, out_s3369, out_e3369, result3369);
PE P3370(out_s3306, out_e3369, clk, rst, out_s3370, out_e3370, result3370);
PE P3371(out_s3307, out_e3370, clk, rst, out_s3371, out_e3371, result3371);
PE P3372(out_s3308, out_e3371, clk, rst, out_s3372, out_e3372, result3372);
PE P3373(out_s3309, out_e3372, clk, rst, out_s3373, out_e3373, result3373);
PE P3374(out_s3310, out_e3373, clk, rst, out_s3374, out_e3374, result3374);
PE P3375(out_s3311, out_e3374, clk, rst, out_s3375, out_e3375, result3375);
PE P3376(out_s3312, out_e3375, clk, rst, out_s3376, out_e3376, result3376);
PE P3377(out_s3313, out_e3376, clk, rst, out_s3377, out_e3377, result3377);
PE P3378(out_s3314, out_e3377, clk, rst, out_s3378, out_e3378, result3378);
PE P3379(out_s3315, out_e3378, clk, rst, out_s3379, out_e3379, result3379);
PE P3380(out_s3316, out_e3379, clk, rst, out_s3380, out_e3380, result3380);
PE P3381(out_s3317, out_e3380, clk, rst, out_s3381, out_e3381, result3381);
PE P3382(out_s3318, out_e3381, clk, rst, out_s3382, out_e3382, result3382);
PE P3383(out_s3319, out_e3382, clk, rst, out_s3383, out_e3383, result3383);
PE P3384(out_s3320, out_e3383, clk, rst, out_s3384, out_e3384, result3384);
PE P3385(out_s3321, out_e3384, clk, rst, out_s3385, out_e3385, result3385);
PE P3386(out_s3322, out_e3385, clk, rst, out_s3386, out_e3386, result3386);
PE P3387(out_s3323, out_e3386, clk, rst, out_s3387, out_e3387, result3387);
PE P3388(out_s3324, out_e3387, clk, rst, out_s3388, out_e3388, result3388);
PE P3389(out_s3325, out_e3388, clk, rst, out_s3389, out_e3389, result3389);
PE P3390(out_s3326, out_e3389, clk, rst, out_s3390, out_e3390, result3390);
PE P3391(out_s3327, out_e3390, clk, rst, out_s3391, out_e3391, result3391);

PE P3393(out_s3329, out_e3392, clk, rst, out_s3393, out_e3393, result3393);
PE P3394(out_s3330, out_e3393, clk, rst, out_s3394, out_e3394, result3394);
PE P3395(out_s3331, out_e3394, clk, rst, out_s3395, out_e3395, result3395);
PE P3396(out_s3332, out_e3395, clk, rst, out_s3396, out_e3396, result3396);
PE P3397(out_s3333, out_e3396, clk, rst, out_s3397, out_e3397, result3397);
PE P3398(out_s3334, out_e3397, clk, rst, out_s3398, out_e3398, result3398);
PE P3399(out_s3335, out_e3398, clk, rst, out_s3399, out_e3399, result3399);
PE P3400(out_s3336, out_e3399, clk, rst, out_s3400, out_e3400, result3400);
PE P3401(out_s3337, out_e3400, clk, rst, out_s3401, out_e3401, result3401);
PE P3402(out_s3338, out_e3401, clk, rst, out_s3402, out_e3402, result3402);
PE P3403(out_s3339, out_e3402, clk, rst, out_s3403, out_e3403, result3403);
PE P3404(out_s3340, out_e3403, clk, rst, out_s3404, out_e3404, result3404);
PE P3405(out_s3341, out_e3404, clk, rst, out_s3405, out_e3405, result3405);
PE P3406(out_s3342, out_e3405, clk, rst, out_s3406, out_e3406, result3406);
PE P3407(out_s3343, out_e3406, clk, rst, out_s3407, out_e3407, result3407);
PE P3408(out_s3344, out_e3407, clk, rst, out_s3408, out_e3408, result3408);
PE P3409(out_s3345, out_e3408, clk, rst, out_s3409, out_e3409, result3409);
PE P3410(out_s3346, out_e3409, clk, rst, out_s3410, out_e3410, result3410);
PE P3411(out_s3347, out_e3410, clk, rst, out_s3411, out_e3411, result3411);
PE P3412(out_s3348, out_e3411, clk, rst, out_s3412, out_e3412, result3412);
PE P3413(out_s3349, out_e3412, clk, rst, out_s3413, out_e3413, result3413);
PE P3414(out_s3350, out_e3413, clk, rst, out_s3414, out_e3414, result3414);
PE P3415(out_s3351, out_e3414, clk, rst, out_s3415, out_e3415, result3415);
PE P3416(out_s3352, out_e3415, clk, rst, out_s3416, out_e3416, result3416);
PE P3417(out_s3353, out_e3416, clk, rst, out_s3417, out_e3417, result3417);
PE P3418(out_s3354, out_e3417, clk, rst, out_s3418, out_e3418, result3418);
PE P3419(out_s3355, out_e3418, clk, rst, out_s3419, out_e3419, result3419);
PE P3420(out_s3356, out_e3419, clk, rst, out_s3420, out_e3420, result3420);
PE P3421(out_s3357, out_e3420, clk, rst, out_s3421, out_e3421, result3421);
PE P3422(out_s3358, out_e3421, clk, rst, out_s3422, out_e3422, result3422);
PE P3423(out_s3359, out_e3422, clk, rst, out_s3423, out_e3423, result3423);
PE P3424(out_s3360, out_e3423, clk, rst, out_s3424, out_e3424, result3424);
PE P3425(out_s3361, out_e3424, clk, rst, out_s3425, out_e3425, result3425);
PE P3426(out_s3362, out_e3425, clk, rst, out_s3426, out_e3426, result3426);
PE P3427(out_s3363, out_e3426, clk, rst, out_s3427, out_e3427, result3427);
PE P3428(out_s3364, out_e3427, clk, rst, out_s3428, out_e3428, result3428);
PE P3429(out_s3365, out_e3428, clk, rst, out_s3429, out_e3429, result3429);
PE P3430(out_s3366, out_e3429, clk, rst, out_s3430, out_e3430, result3430);
PE P3431(out_s3367, out_e3430, clk, rst, out_s3431, out_e3431, result3431);
PE P3432(out_s3368, out_e3431, clk, rst, out_s3432, out_e3432, result3432);
PE P3433(out_s3369, out_e3432, clk, rst, out_s3433, out_e3433, result3433);
PE P3434(out_s3370, out_e3433, clk, rst, out_s3434, out_e3434, result3434);
PE P3435(out_s3371, out_e3434, clk, rst, out_s3435, out_e3435, result3435);
PE P3436(out_s3372, out_e3435, clk, rst, out_s3436, out_e3436, result3436);
PE P3437(out_s3373, out_e3436, clk, rst, out_s3437, out_e3437, result3437);
PE P3438(out_s3374, out_e3437, clk, rst, out_s3438, out_e3438, result3438);
PE P3439(out_s3375, out_e3438, clk, rst, out_s3439, out_e3439, result3439);
PE P3440(out_s3376, out_e3439, clk, rst, out_s3440, out_e3440, result3440);
PE P3441(out_s3377, out_e3440, clk, rst, out_s3441, out_e3441, result3441);
PE P3442(out_s3378, out_e3441, clk, rst, out_s3442, out_e3442, result3442);
PE P3443(out_s3379, out_e3442, clk, rst, out_s3443, out_e3443, result3443);
PE P3444(out_s3380, out_e3443, clk, rst, out_s3444, out_e3444, result3444);
PE P3445(out_s3381, out_e3444, clk, rst, out_s3445, out_e3445, result3445);
PE P3446(out_s3382, out_e3445, clk, rst, out_s3446, out_e3446, result3446);
PE P3447(out_s3383, out_e3446, clk, rst, out_s3447, out_e3447, result3447);
PE P3448(out_s3384, out_e3447, clk, rst, out_s3448, out_e3448, result3448);
PE P3449(out_s3385, out_e3448, clk, rst, out_s3449, out_e3449, result3449);
PE P3450(out_s3386, out_e3449, clk, rst, out_s3450, out_e3450, result3450);
PE P3451(out_s3387, out_e3450, clk, rst, out_s3451, out_e3451, result3451);
PE P3452(out_s3388, out_e3451, clk, rst, out_s3452, out_e3452, result3452);
PE P3453(out_s3389, out_e3452, clk, rst, out_s3453, out_e3453, result3453);
PE P3454(out_s3390, out_e3453, clk, rst, out_s3454, out_e3454, result3454);
PE P3455(out_s3391, out_e3454, clk, rst, out_s3455, out_e3455, result3455);

PE P3457(out_s3393, out_e3456, clk, rst, out_s3457, out_e3457, result3457);
PE P3458(out_s3394, out_e3457, clk, rst, out_s3458, out_e3458, result3458);
PE P3459(out_s3395, out_e3458, clk, rst, out_s3459, out_e3459, result3459);
PE P3460(out_s3396, out_e3459, clk, rst, out_s3460, out_e3460, result3460);
PE P3461(out_s3397, out_e3460, clk, rst, out_s3461, out_e3461, result3461);
PE P3462(out_s3398, out_e3461, clk, rst, out_s3462, out_e3462, result3462);
PE P3463(out_s3399, out_e3462, clk, rst, out_s3463, out_e3463, result3463);
PE P3464(out_s3400, out_e3463, clk, rst, out_s3464, out_e3464, result3464);
PE P3465(out_s3401, out_e3464, clk, rst, out_s3465, out_e3465, result3465);
PE P3466(out_s3402, out_e3465, clk, rst, out_s3466, out_e3466, result3466);
PE P3467(out_s3403, out_e3466, clk, rst, out_s3467, out_e3467, result3467);
PE P3468(out_s3404, out_e3467, clk, rst, out_s3468, out_e3468, result3468);
PE P3469(out_s3405, out_e3468, clk, rst, out_s3469, out_e3469, result3469);
PE P3470(out_s3406, out_e3469, clk, rst, out_s3470, out_e3470, result3470);
PE P3471(out_s3407, out_e3470, clk, rst, out_s3471, out_e3471, result3471);
PE P3472(out_s3408, out_e3471, clk, rst, out_s3472, out_e3472, result3472);
PE P3473(out_s3409, out_e3472, clk, rst, out_s3473, out_e3473, result3473);
PE P3474(out_s3410, out_e3473, clk, rst, out_s3474, out_e3474, result3474);
PE P3475(out_s3411, out_e3474, clk, rst, out_s3475, out_e3475, result3475);
PE P3476(out_s3412, out_e3475, clk, rst, out_s3476, out_e3476, result3476);
PE P3477(out_s3413, out_e3476, clk, rst, out_s3477, out_e3477, result3477);
PE P3478(out_s3414, out_e3477, clk, rst, out_s3478, out_e3478, result3478);
PE P3479(out_s3415, out_e3478, clk, rst, out_s3479, out_e3479, result3479);
PE P3480(out_s3416, out_e3479, clk, rst, out_s3480, out_e3480, result3480);
PE P3481(out_s3417, out_e3480, clk, rst, out_s3481, out_e3481, result3481);
PE P3482(out_s3418, out_e3481, clk, rst, out_s3482, out_e3482, result3482);
PE P3483(out_s3419, out_e3482, clk, rst, out_s3483, out_e3483, result3483);
PE P3484(out_s3420, out_e3483, clk, rst, out_s3484, out_e3484, result3484);
PE P3485(out_s3421, out_e3484, clk, rst, out_s3485, out_e3485, result3485);
PE P3486(out_s3422, out_e3485, clk, rst, out_s3486, out_e3486, result3486);
PE P3487(out_s3423, out_e3486, clk, rst, out_s3487, out_e3487, result3487);
PE P3488(out_s3424, out_e3487, clk, rst, out_s3488, out_e3488, result3488);
PE P3489(out_s3425, out_e3488, clk, rst, out_s3489, out_e3489, result3489);
PE P3490(out_s3426, out_e3489, clk, rst, out_s3490, out_e3490, result3490);
PE P3491(out_s3427, out_e3490, clk, rst, out_s3491, out_e3491, result3491);
PE P3492(out_s3428, out_e3491, clk, rst, out_s3492, out_e3492, result3492);
PE P3493(out_s3429, out_e3492, clk, rst, out_s3493, out_e3493, result3493);
PE P3494(out_s3430, out_e3493, clk, rst, out_s3494, out_e3494, result3494);
PE P3495(out_s3431, out_e3494, clk, rst, out_s3495, out_e3495, result3495);
PE P3496(out_s3432, out_e3495, clk, rst, out_s3496, out_e3496, result3496);
PE P3497(out_s3433, out_e3496, clk, rst, out_s3497, out_e3497, result3497);
PE P3498(out_s3434, out_e3497, clk, rst, out_s3498, out_e3498, result3498);
PE P3499(out_s3435, out_e3498, clk, rst, out_s3499, out_e3499, result3499);
PE P3500(out_s3436, out_e3499, clk, rst, out_s3500, out_e3500, result3500);
PE P3501(out_s3437, out_e3500, clk, rst, out_s3501, out_e3501, result3501);
PE P3502(out_s3438, out_e3501, clk, rst, out_s3502, out_e3502, result3502);
PE P3503(out_s3439, out_e3502, clk, rst, out_s3503, out_e3503, result3503);
PE P3504(out_s3440, out_e3503, clk, rst, out_s3504, out_e3504, result3504);
PE P3505(out_s3441, out_e3504, clk, rst, out_s3505, out_e3505, result3505);
PE P3506(out_s3442, out_e3505, clk, rst, out_s3506, out_e3506, result3506);
PE P3507(out_s3443, out_e3506, clk, rst, out_s3507, out_e3507, result3507);
PE P3508(out_s3444, out_e3507, clk, rst, out_s3508, out_e3508, result3508);
PE P3509(out_s3445, out_e3508, clk, rst, out_s3509, out_e3509, result3509);
PE P3510(out_s3446, out_e3509, clk, rst, out_s3510, out_e3510, result3510);
PE P3511(out_s3447, out_e3510, clk, rst, out_s3511, out_e3511, result3511);
PE P3512(out_s3448, out_e3511, clk, rst, out_s3512, out_e3512, result3512);
PE P3513(out_s3449, out_e3512, clk, rst, out_s3513, out_e3513, result3513);
PE P3514(out_s3450, out_e3513, clk, rst, out_s3514, out_e3514, result3514);
PE P3515(out_s3451, out_e3514, clk, rst, out_s3515, out_e3515, result3515);
PE P3516(out_s3452, out_e3515, clk, rst, out_s3516, out_e3516, result3516);
PE P3517(out_s3453, out_e3516, clk, rst, out_s3517, out_e3517, result3517);
PE P3518(out_s3454, out_e3517, clk, rst, out_s3518, out_e3518, result3518);
PE P3519(out_s3455, out_e3518, clk, rst, out_s3519, out_e3519, result3519);

PE P3521(out_s3457, out_e3520, clk, rst, out_s3521, out_e3521, result3521);
PE P3522(out_s3458, out_e3521, clk, rst, out_s3522, out_e3522, result3522);
PE P3523(out_s3459, out_e3522, clk, rst, out_s3523, out_e3523, result3523);
PE P3524(out_s3460, out_e3523, clk, rst, out_s3524, out_e3524, result3524);
PE P3525(out_s3461, out_e3524, clk, rst, out_s3525, out_e3525, result3525);
PE P3526(out_s3462, out_e3525, clk, rst, out_s3526, out_e3526, result3526);
PE P3527(out_s3463, out_e3526, clk, rst, out_s3527, out_e3527, result3527);
PE P3528(out_s3464, out_e3527, clk, rst, out_s3528, out_e3528, result3528);
PE P3529(out_s3465, out_e3528, clk, rst, out_s3529, out_e3529, result3529);
PE P3530(out_s3466, out_e3529, clk, rst, out_s3530, out_e3530, result3530);
PE P3531(out_s3467, out_e3530, clk, rst, out_s3531, out_e3531, result3531);
PE P3532(out_s3468, out_e3531, clk, rst, out_s3532, out_e3532, result3532);
PE P3533(out_s3469, out_e3532, clk, rst, out_s3533, out_e3533, result3533);
PE P3534(out_s3470, out_e3533, clk, rst, out_s3534, out_e3534, result3534);
PE P3535(out_s3471, out_e3534, clk, rst, out_s3535, out_e3535, result3535);
PE P3536(out_s3472, out_e3535, clk, rst, out_s3536, out_e3536, result3536);
PE P3537(out_s3473, out_e3536, clk, rst, out_s3537, out_e3537, result3537);
PE P3538(out_s3474, out_e3537, clk, rst, out_s3538, out_e3538, result3538);
PE P3539(out_s3475, out_e3538, clk, rst, out_s3539, out_e3539, result3539);
PE P3540(out_s3476, out_e3539, clk, rst, out_s3540, out_e3540, result3540);
PE P3541(out_s3477, out_e3540, clk, rst, out_s3541, out_e3541, result3541);
PE P3542(out_s3478, out_e3541, clk, rst, out_s3542, out_e3542, result3542);
PE P3543(out_s3479, out_e3542, clk, rst, out_s3543, out_e3543, result3543);
PE P3544(out_s3480, out_e3543, clk, rst, out_s3544, out_e3544, result3544);
PE P3545(out_s3481, out_e3544, clk, rst, out_s3545, out_e3545, result3545);
PE P3546(out_s3482, out_e3545, clk, rst, out_s3546, out_e3546, result3546);
PE P3547(out_s3483, out_e3546, clk, rst, out_s3547, out_e3547, result3547);
PE P3548(out_s3484, out_e3547, clk, rst, out_s3548, out_e3548, result3548);
PE P3549(out_s3485, out_e3548, clk, rst, out_s3549, out_e3549, result3549);
PE P3550(out_s3486, out_e3549, clk, rst, out_s3550, out_e3550, result3550);
PE P3551(out_s3487, out_e3550, clk, rst, out_s3551, out_e3551, result3551);
PE P3552(out_s3488, out_e3551, clk, rst, out_s3552, out_e3552, result3552);
PE P3553(out_s3489, out_e3552, clk, rst, out_s3553, out_e3553, result3553);
PE P3554(out_s3490, out_e3553, clk, rst, out_s3554, out_e3554, result3554);
PE P3555(out_s3491, out_e3554, clk, rst, out_s3555, out_e3555, result3555);
PE P3556(out_s3492, out_e3555, clk, rst, out_s3556, out_e3556, result3556);
PE P3557(out_s3493, out_e3556, clk, rst, out_s3557, out_e3557, result3557);
PE P3558(out_s3494, out_e3557, clk, rst, out_s3558, out_e3558, result3558);
PE P3559(out_s3495, out_e3558, clk, rst, out_s3559, out_e3559, result3559);
PE P3560(out_s3496, out_e3559, clk, rst, out_s3560, out_e3560, result3560);
PE P3561(out_s3497, out_e3560, clk, rst, out_s3561, out_e3561, result3561);
PE P3562(out_s3498, out_e3561, clk, rst, out_s3562, out_e3562, result3562);
PE P3563(out_s3499, out_e3562, clk, rst, out_s3563, out_e3563, result3563);
PE P3564(out_s3500, out_e3563, clk, rst, out_s3564, out_e3564, result3564);
PE P3565(out_s3501, out_e3564, clk, rst, out_s3565, out_e3565, result3565);
PE P3566(out_s3502, out_e3565, clk, rst, out_s3566, out_e3566, result3566);
PE P3567(out_s3503, out_e3566, clk, rst, out_s3567, out_e3567, result3567);
PE P3568(out_s3504, out_e3567, clk, rst, out_s3568, out_e3568, result3568);
PE P3569(out_s3505, out_e3568, clk, rst, out_s3569, out_e3569, result3569);
PE P3570(out_s3506, out_e3569, clk, rst, out_s3570, out_e3570, result3570);
PE P3571(out_s3507, out_e3570, clk, rst, out_s3571, out_e3571, result3571);
PE P3572(out_s3508, out_e3571, clk, rst, out_s3572, out_e3572, result3572);
PE P3573(out_s3509, out_e3572, clk, rst, out_s3573, out_e3573, result3573);
PE P3574(out_s3510, out_e3573, clk, rst, out_s3574, out_e3574, result3574);
PE P3575(out_s3511, out_e3574, clk, rst, out_s3575, out_e3575, result3575);
PE P3576(out_s3512, out_e3575, clk, rst, out_s3576, out_e3576, result3576);
PE P3577(out_s3513, out_e3576, clk, rst, out_s3577, out_e3577, result3577);
PE P3578(out_s3514, out_e3577, clk, rst, out_s3578, out_e3578, result3578);
PE P3579(out_s3515, out_e3578, clk, rst, out_s3579, out_e3579, result3579);
PE P3580(out_s3516, out_e3579, clk, rst, out_s3580, out_e3580, result3580);
PE P3581(out_s3517, out_e3580, clk, rst, out_s3581, out_e3581, result3581);
PE P3582(out_s3518, out_e3581, clk, rst, out_s3582, out_e3582, result3582);
PE P3583(out_s3519, out_e3582, clk, rst, out_s3583, out_e3583, result3583);

PE P3585(out_s3521, out_e3584, clk, rst, out_s3585, out_e3585, result3585);
PE P3586(out_s3522, out_e3585, clk, rst, out_s3586, out_e3586, result3586);
PE P3587(out_s3523, out_e3586, clk, rst, out_s3587, out_e3587, result3587);
PE P3588(out_s3524, out_e3587, clk, rst, out_s3588, out_e3588, result3588);
PE P3589(out_s3525, out_e3588, clk, rst, out_s3589, out_e3589, result3589);
PE P3590(out_s3526, out_e3589, clk, rst, out_s3590, out_e3590, result3590);
PE P3591(out_s3527, out_e3590, clk, rst, out_s3591, out_e3591, result3591);
PE P3592(out_s3528, out_e3591, clk, rst, out_s3592, out_e3592, result3592);
PE P3593(out_s3529, out_e3592, clk, rst, out_s3593, out_e3593, result3593);
PE P3594(out_s3530, out_e3593, clk, rst, out_s3594, out_e3594, result3594);
PE P3595(out_s3531, out_e3594, clk, rst, out_s3595, out_e3595, result3595);
PE P3596(out_s3532, out_e3595, clk, rst, out_s3596, out_e3596, result3596);
PE P3597(out_s3533, out_e3596, clk, rst, out_s3597, out_e3597, result3597);
PE P3598(out_s3534, out_e3597, clk, rst, out_s3598, out_e3598, result3598);
PE P3599(out_s3535, out_e3598, clk, rst, out_s3599, out_e3599, result3599);
PE P3600(out_s3536, out_e3599, clk, rst, out_s3600, out_e3600, result3600);
PE P3601(out_s3537, out_e3600, clk, rst, out_s3601, out_e3601, result3601);
PE P3602(out_s3538, out_e3601, clk, rst, out_s3602, out_e3602, result3602);
PE P3603(out_s3539, out_e3602, clk, rst, out_s3603, out_e3603, result3603);
PE P3604(out_s3540, out_e3603, clk, rst, out_s3604, out_e3604, result3604);
PE P3605(out_s3541, out_e3604, clk, rst, out_s3605, out_e3605, result3605);
PE P3606(out_s3542, out_e3605, clk, rst, out_s3606, out_e3606, result3606);
PE P3607(out_s3543, out_e3606, clk, rst, out_s3607, out_e3607, result3607);
PE P3608(out_s3544, out_e3607, clk, rst, out_s3608, out_e3608, result3608);
PE P3609(out_s3545, out_e3608, clk, rst, out_s3609, out_e3609, result3609);
PE P3610(out_s3546, out_e3609, clk, rst, out_s3610, out_e3610, result3610);
PE P3611(out_s3547, out_e3610, clk, rst, out_s3611, out_e3611, result3611);
PE P3612(out_s3548, out_e3611, clk, rst, out_s3612, out_e3612, result3612);
PE P3613(out_s3549, out_e3612, clk, rst, out_s3613, out_e3613, result3613);
PE P3614(out_s3550, out_e3613, clk, rst, out_s3614, out_e3614, result3614);
PE P3615(out_s3551, out_e3614, clk, rst, out_s3615, out_e3615, result3615);
PE P3616(out_s3552, out_e3615, clk, rst, out_s3616, out_e3616, result3616);
PE P3617(out_s3553, out_e3616, clk, rst, out_s3617, out_e3617, result3617);
PE P3618(out_s3554, out_e3617, clk, rst, out_s3618, out_e3618, result3618);
PE P3619(out_s3555, out_e3618, clk, rst, out_s3619, out_e3619, result3619);
PE P3620(out_s3556, out_e3619, clk, rst, out_s3620, out_e3620, result3620);
PE P3621(out_s3557, out_e3620, clk, rst, out_s3621, out_e3621, result3621);
PE P3622(out_s3558, out_e3621, clk, rst, out_s3622, out_e3622, result3622);
PE P3623(out_s3559, out_e3622, clk, rst, out_s3623, out_e3623, result3623);
PE P3624(out_s3560, out_e3623, clk, rst, out_s3624, out_e3624, result3624);
PE P3625(out_s3561, out_e3624, clk, rst, out_s3625, out_e3625, result3625);
PE P3626(out_s3562, out_e3625, clk, rst, out_s3626, out_e3626, result3626);
PE P3627(out_s3563, out_e3626, clk, rst, out_s3627, out_e3627, result3627);
PE P3628(out_s3564, out_e3627, clk, rst, out_s3628, out_e3628, result3628);
PE P3629(out_s3565, out_e3628, clk, rst, out_s3629, out_e3629, result3629);
PE P3630(out_s3566, out_e3629, clk, rst, out_s3630, out_e3630, result3630);
PE P3631(out_s3567, out_e3630, clk, rst, out_s3631, out_e3631, result3631);
PE P3632(out_s3568, out_e3631, clk, rst, out_s3632, out_e3632, result3632);
PE P3633(out_s3569, out_e3632, clk, rst, out_s3633, out_e3633, result3633);
PE P3634(out_s3570, out_e3633, clk, rst, out_s3634, out_e3634, result3634);
PE P3635(out_s3571, out_e3634, clk, rst, out_s3635, out_e3635, result3635);
PE P3636(out_s3572, out_e3635, clk, rst, out_s3636, out_e3636, result3636);
PE P3637(out_s3573, out_e3636, clk, rst, out_s3637, out_e3637, result3637);
PE P3638(out_s3574, out_e3637, clk, rst, out_s3638, out_e3638, result3638);
PE P3639(out_s3575, out_e3638, clk, rst, out_s3639, out_e3639, result3639);
PE P3640(out_s3576, out_e3639, clk, rst, out_s3640, out_e3640, result3640);
PE P3641(out_s3577, out_e3640, clk, rst, out_s3641, out_e3641, result3641);
PE P3642(out_s3578, out_e3641, clk, rst, out_s3642, out_e3642, result3642);
PE P3643(out_s3579, out_e3642, clk, rst, out_s3643, out_e3643, result3643);
PE P3644(out_s3580, out_e3643, clk, rst, out_s3644, out_e3644, result3644);
PE P3645(out_s3581, out_e3644, clk, rst, out_s3645, out_e3645, result3645);
PE P3646(out_s3582, out_e3645, clk, rst, out_s3646, out_e3646, result3646);
PE P3647(out_s3583, out_e3646, clk, rst, out_s3647, out_e3647, result3647);

PE P3649(out_s3585, out_e3648, clk, rst, out_s3649, out_e3649, result3649);
PE P3650(out_s3586, out_e3649, clk, rst, out_s3650, out_e3650, result3650);
PE P3651(out_s3587, out_e3650, clk, rst, out_s3651, out_e3651, result3651);
PE P3652(out_s3588, out_e3651, clk, rst, out_s3652, out_e3652, result3652);
PE P3653(out_s3589, out_e3652, clk, rst, out_s3653, out_e3653, result3653);
PE P3654(out_s3590, out_e3653, clk, rst, out_s3654, out_e3654, result3654);
PE P3655(out_s3591, out_e3654, clk, rst, out_s3655, out_e3655, result3655);
PE P3656(out_s3592, out_e3655, clk, rst, out_s3656, out_e3656, result3656);
PE P3657(out_s3593, out_e3656, clk, rst, out_s3657, out_e3657, result3657);
PE P3658(out_s3594, out_e3657, clk, rst, out_s3658, out_e3658, result3658);
PE P3659(out_s3595, out_e3658, clk, rst, out_s3659, out_e3659, result3659);
PE P3660(out_s3596, out_e3659, clk, rst, out_s3660, out_e3660, result3660);
PE P3661(out_s3597, out_e3660, clk, rst, out_s3661, out_e3661, result3661);
PE P3662(out_s3598, out_e3661, clk, rst, out_s3662, out_e3662, result3662);
PE P3663(out_s3599, out_e3662, clk, rst, out_s3663, out_e3663, result3663);
PE P3664(out_s3600, out_e3663, clk, rst, out_s3664, out_e3664, result3664);
PE P3665(out_s3601, out_e3664, clk, rst, out_s3665, out_e3665, result3665);
PE P3666(out_s3602, out_e3665, clk, rst, out_s3666, out_e3666, result3666);
PE P3667(out_s3603, out_e3666, clk, rst, out_s3667, out_e3667, result3667);
PE P3668(out_s3604, out_e3667, clk, rst, out_s3668, out_e3668, result3668);
PE P3669(out_s3605, out_e3668, clk, rst, out_s3669, out_e3669, result3669);
PE P3670(out_s3606, out_e3669, clk, rst, out_s3670, out_e3670, result3670);
PE P3671(out_s3607, out_e3670, clk, rst, out_s3671, out_e3671, result3671);
PE P3672(out_s3608, out_e3671, clk, rst, out_s3672, out_e3672, result3672);
PE P3673(out_s3609, out_e3672, clk, rst, out_s3673, out_e3673, result3673);
PE P3674(out_s3610, out_e3673, clk, rst, out_s3674, out_e3674, result3674);
PE P3675(out_s3611, out_e3674, clk, rst, out_s3675, out_e3675, result3675);
PE P3676(out_s3612, out_e3675, clk, rst, out_s3676, out_e3676, result3676);
PE P3677(out_s3613, out_e3676, clk, rst, out_s3677, out_e3677, result3677);
PE P3678(out_s3614, out_e3677, clk, rst, out_s3678, out_e3678, result3678);
PE P3679(out_s3615, out_e3678, clk, rst, out_s3679, out_e3679, result3679);
PE P3680(out_s3616, out_e3679, clk, rst, out_s3680, out_e3680, result3680);
PE P3681(out_s3617, out_e3680, clk, rst, out_s3681, out_e3681, result3681);
PE P3682(out_s3618, out_e3681, clk, rst, out_s3682, out_e3682, result3682);
PE P3683(out_s3619, out_e3682, clk, rst, out_s3683, out_e3683, result3683);
PE P3684(out_s3620, out_e3683, clk, rst, out_s3684, out_e3684, result3684);
PE P3685(out_s3621, out_e3684, clk, rst, out_s3685, out_e3685, result3685);
PE P3686(out_s3622, out_e3685, clk, rst, out_s3686, out_e3686, result3686);
PE P3687(out_s3623, out_e3686, clk, rst, out_s3687, out_e3687, result3687);
PE P3688(out_s3624, out_e3687, clk, rst, out_s3688, out_e3688, result3688);
PE P3689(out_s3625, out_e3688, clk, rst, out_s3689, out_e3689, result3689);
PE P3690(out_s3626, out_e3689, clk, rst, out_s3690, out_e3690, result3690);
PE P3691(out_s3627, out_e3690, clk, rst, out_s3691, out_e3691, result3691);
PE P3692(out_s3628, out_e3691, clk, rst, out_s3692, out_e3692, result3692);
PE P3693(out_s3629, out_e3692, clk, rst, out_s3693, out_e3693, result3693);
PE P3694(out_s3630, out_e3693, clk, rst, out_s3694, out_e3694, result3694);
PE P3695(out_s3631, out_e3694, clk, rst, out_s3695, out_e3695, result3695);
PE P3696(out_s3632, out_e3695, clk, rst, out_s3696, out_e3696, result3696);
PE P3697(out_s3633, out_e3696, clk, rst, out_s3697, out_e3697, result3697);
PE P3698(out_s3634, out_e3697, clk, rst, out_s3698, out_e3698, result3698);
PE P3699(out_s3635, out_e3698, clk, rst, out_s3699, out_e3699, result3699);
PE P3700(out_s3636, out_e3699, clk, rst, out_s3700, out_e3700, result3700);
PE P3701(out_s3637, out_e3700, clk, rst, out_s3701, out_e3701, result3701);
PE P3702(out_s3638, out_e3701, clk, rst, out_s3702, out_e3702, result3702);
PE P3703(out_s3639, out_e3702, clk, rst, out_s3703, out_e3703, result3703);
PE P3704(out_s3640, out_e3703, clk, rst, out_s3704, out_e3704, result3704);
PE P3705(out_s3641, out_e3704, clk, rst, out_s3705, out_e3705, result3705);
PE P3706(out_s3642, out_e3705, clk, rst, out_s3706, out_e3706, result3706);
PE P3707(out_s3643, out_e3706, clk, rst, out_s3707, out_e3707, result3707);
PE P3708(out_s3644, out_e3707, clk, rst, out_s3708, out_e3708, result3708);
PE P3709(out_s3645, out_e3708, clk, rst, out_s3709, out_e3709, result3709);
PE P3710(out_s3646, out_e3709, clk, rst, out_s3710, out_e3710, result3710);
PE P3711(out_s3647, out_e3710, clk, rst, out_s3711, out_e3711, result3711);

PE P3713(out_s3649, out_e3712, clk, rst, out_s3713, out_e3713, result3713);
PE P3714(out_s3650, out_e3713, clk, rst, out_s3714, out_e3714, result3714);
PE P3715(out_s3651, out_e3714, clk, rst, out_s3715, out_e3715, result3715);
PE P3716(out_s3652, out_e3715, clk, rst, out_s3716, out_e3716, result3716);
PE P3717(out_s3653, out_e3716, clk, rst, out_s3717, out_e3717, result3717);
PE P3718(out_s3654, out_e3717, clk, rst, out_s3718, out_e3718, result3718);
PE P3719(out_s3655, out_e3718, clk, rst, out_s3719, out_e3719, result3719);
PE P3720(out_s3656, out_e3719, clk, rst, out_s3720, out_e3720, result3720);
PE P3721(out_s3657, out_e3720, clk, rst, out_s3721, out_e3721, result3721);
PE P3722(out_s3658, out_e3721, clk, rst, out_s3722, out_e3722, result3722);
PE P3723(out_s3659, out_e3722, clk, rst, out_s3723, out_e3723, result3723);
PE P3724(out_s3660, out_e3723, clk, rst, out_s3724, out_e3724, result3724);
PE P3725(out_s3661, out_e3724, clk, rst, out_s3725, out_e3725, result3725);
PE P3726(out_s3662, out_e3725, clk, rst, out_s3726, out_e3726, result3726);
PE P3727(out_s3663, out_e3726, clk, rst, out_s3727, out_e3727, result3727);
PE P3728(out_s3664, out_e3727, clk, rst, out_s3728, out_e3728, result3728);
PE P3729(out_s3665, out_e3728, clk, rst, out_s3729, out_e3729, result3729);
PE P3730(out_s3666, out_e3729, clk, rst, out_s3730, out_e3730, result3730);
PE P3731(out_s3667, out_e3730, clk, rst, out_s3731, out_e3731, result3731);
PE P3732(out_s3668, out_e3731, clk, rst, out_s3732, out_e3732, result3732);
PE P3733(out_s3669, out_e3732, clk, rst, out_s3733, out_e3733, result3733);
PE P3734(out_s3670, out_e3733, clk, rst, out_s3734, out_e3734, result3734);
PE P3735(out_s3671, out_e3734, clk, rst, out_s3735, out_e3735, result3735);
PE P3736(out_s3672, out_e3735, clk, rst, out_s3736, out_e3736, result3736);
PE P3737(out_s3673, out_e3736, clk, rst, out_s3737, out_e3737, result3737);
PE P3738(out_s3674, out_e3737, clk, rst, out_s3738, out_e3738, result3738);
PE P3739(out_s3675, out_e3738, clk, rst, out_s3739, out_e3739, result3739);
PE P3740(out_s3676, out_e3739, clk, rst, out_s3740, out_e3740, result3740);
PE P3741(out_s3677, out_e3740, clk, rst, out_s3741, out_e3741, result3741);
PE P3742(out_s3678, out_e3741, clk, rst, out_s3742, out_e3742, result3742);
PE P3743(out_s3679, out_e3742, clk, rst, out_s3743, out_e3743, result3743);
PE P3744(out_s3680, out_e3743, clk, rst, out_s3744, out_e3744, result3744);
PE P3745(out_s3681, out_e3744, clk, rst, out_s3745, out_e3745, result3745);
PE P3746(out_s3682, out_e3745, clk, rst, out_s3746, out_e3746, result3746);
PE P3747(out_s3683, out_e3746, clk, rst, out_s3747, out_e3747, result3747);
PE P3748(out_s3684, out_e3747, clk, rst, out_s3748, out_e3748, result3748);
PE P3749(out_s3685, out_e3748, clk, rst, out_s3749, out_e3749, result3749);
PE P3750(out_s3686, out_e3749, clk, rst, out_s3750, out_e3750, result3750);
PE P3751(out_s3687, out_e3750, clk, rst, out_s3751, out_e3751, result3751);
PE P3752(out_s3688, out_e3751, clk, rst, out_s3752, out_e3752, result3752);
PE P3753(out_s3689, out_e3752, clk, rst, out_s3753, out_e3753, result3753);
PE P3754(out_s3690, out_e3753, clk, rst, out_s3754, out_e3754, result3754);
PE P3755(out_s3691, out_e3754, clk, rst, out_s3755, out_e3755, result3755);
PE P3756(out_s3692, out_e3755, clk, rst, out_s3756, out_e3756, result3756);
PE P3757(out_s3693, out_e3756, clk, rst, out_s3757, out_e3757, result3757);
PE P3758(out_s3694, out_e3757, clk, rst, out_s3758, out_e3758, result3758);
PE P3759(out_s3695, out_e3758, clk, rst, out_s3759, out_e3759, result3759);
PE P3760(out_s3696, out_e3759, clk, rst, out_s3760, out_e3760, result3760);
PE P3761(out_s3697, out_e3760, clk, rst, out_s3761, out_e3761, result3761);
PE P3762(out_s3698, out_e3761, clk, rst, out_s3762, out_e3762, result3762);
PE P3763(out_s3699, out_e3762, clk, rst, out_s3763, out_e3763, result3763);
PE P3764(out_s3700, out_e3763, clk, rst, out_s3764, out_e3764, result3764);
PE P3765(out_s3701, out_e3764, clk, rst, out_s3765, out_e3765, result3765);
PE P3766(out_s3702, out_e3765, clk, rst, out_s3766, out_e3766, result3766);
PE P3767(out_s3703, out_e3766, clk, rst, out_s3767, out_e3767, result3767);
PE P3768(out_s3704, out_e3767, clk, rst, out_s3768, out_e3768, result3768);
PE P3769(out_s3705, out_e3768, clk, rst, out_s3769, out_e3769, result3769);
PE P3770(out_s3706, out_e3769, clk, rst, out_s3770, out_e3770, result3770);
PE P3771(out_s3707, out_e3770, clk, rst, out_s3771, out_e3771, result3771);
PE P3772(out_s3708, out_e3771, clk, rst, out_s3772, out_e3772, result3772);
PE P3773(out_s3709, out_e3772, clk, rst, out_s3773, out_e3773, result3773);
PE P3774(out_s3710, out_e3773, clk, rst, out_s3774, out_e3774, result3774);
PE P3775(out_s3711, out_e3774, clk, rst, out_s3775, out_e3775, result3775);

PE P3777(out_s3713, out_e3776, clk, rst, out_s3777, out_e3777, result3777);
PE P3778(out_s3714, out_e3777, clk, rst, out_s3778, out_e3778, result3778);
PE P3779(out_s3715, out_e3778, clk, rst, out_s3779, out_e3779, result3779);
PE P3780(out_s3716, out_e3779, clk, rst, out_s3780, out_e3780, result3780);
PE P3781(out_s3717, out_e3780, clk, rst, out_s3781, out_e3781, result3781);
PE P3782(out_s3718, out_e3781, clk, rst, out_s3782, out_e3782, result3782);
PE P3783(out_s3719, out_e3782, clk, rst, out_s3783, out_e3783, result3783);
PE P3784(out_s3720, out_e3783, clk, rst, out_s3784, out_e3784, result3784);
PE P3785(out_s3721, out_e3784, clk, rst, out_s3785, out_e3785, result3785);
PE P3786(out_s3722, out_e3785, clk, rst, out_s3786, out_e3786, result3786);
PE P3787(out_s3723, out_e3786, clk, rst, out_s3787, out_e3787, result3787);
PE P3788(out_s3724, out_e3787, clk, rst, out_s3788, out_e3788, result3788);
PE P3789(out_s3725, out_e3788, clk, rst, out_s3789, out_e3789, result3789);
PE P3790(out_s3726, out_e3789, clk, rst, out_s3790, out_e3790, result3790);
PE P3791(out_s3727, out_e3790, clk, rst, out_s3791, out_e3791, result3791);
PE P3792(out_s3728, out_e3791, clk, rst, out_s3792, out_e3792, result3792);
PE P3793(out_s3729, out_e3792, clk, rst, out_s3793, out_e3793, result3793);
PE P3794(out_s3730, out_e3793, clk, rst, out_s3794, out_e3794, result3794);
PE P3795(out_s3731, out_e3794, clk, rst, out_s3795, out_e3795, result3795);
PE P3796(out_s3732, out_e3795, clk, rst, out_s3796, out_e3796, result3796);
PE P3797(out_s3733, out_e3796, clk, rst, out_s3797, out_e3797, result3797);
PE P3798(out_s3734, out_e3797, clk, rst, out_s3798, out_e3798, result3798);
PE P3799(out_s3735, out_e3798, clk, rst, out_s3799, out_e3799, result3799);
PE P3800(out_s3736, out_e3799, clk, rst, out_s3800, out_e3800, result3800);
PE P3801(out_s3737, out_e3800, clk, rst, out_s3801, out_e3801, result3801);
PE P3802(out_s3738, out_e3801, clk, rst, out_s3802, out_e3802, result3802);
PE P3803(out_s3739, out_e3802, clk, rst, out_s3803, out_e3803, result3803);
PE P3804(out_s3740, out_e3803, clk, rst, out_s3804, out_e3804, result3804);
PE P3805(out_s3741, out_e3804, clk, rst, out_s3805, out_e3805, result3805);
PE P3806(out_s3742, out_e3805, clk, rst, out_s3806, out_e3806, result3806);
PE P3807(out_s3743, out_e3806, clk, rst, out_s3807, out_e3807, result3807);
PE P3808(out_s3744, out_e3807, clk, rst, out_s3808, out_e3808, result3808);
PE P3809(out_s3745, out_e3808, clk, rst, out_s3809, out_e3809, result3809);
PE P3810(out_s3746, out_e3809, clk, rst, out_s3810, out_e3810, result3810);
PE P3811(out_s3747, out_e3810, clk, rst, out_s3811, out_e3811, result3811);
PE P3812(out_s3748, out_e3811, clk, rst, out_s3812, out_e3812, result3812);
PE P3813(out_s3749, out_e3812, clk, rst, out_s3813, out_e3813, result3813);
PE P3814(out_s3750, out_e3813, clk, rst, out_s3814, out_e3814, result3814);
PE P3815(out_s3751, out_e3814, clk, rst, out_s3815, out_e3815, result3815);
PE P3816(out_s3752, out_e3815, clk, rst, out_s3816, out_e3816, result3816);
PE P3817(out_s3753, out_e3816, clk, rst, out_s3817, out_e3817, result3817);
PE P3818(out_s3754, out_e3817, clk, rst, out_s3818, out_e3818, result3818);
PE P3819(out_s3755, out_e3818, clk, rst, out_s3819, out_e3819, result3819);
PE P3820(out_s3756, out_e3819, clk, rst, out_s3820, out_e3820, result3820);
PE P3821(out_s3757, out_e3820, clk, rst, out_s3821, out_e3821, result3821);
PE P3822(out_s3758, out_e3821, clk, rst, out_s3822, out_e3822, result3822);
PE P3823(out_s3759, out_e3822, clk, rst, out_s3823, out_e3823, result3823);
PE P3824(out_s3760, out_e3823, clk, rst, out_s3824, out_e3824, result3824);
PE P3825(out_s3761, out_e3824, clk, rst, out_s3825, out_e3825, result3825);
PE P3826(out_s3762, out_e3825, clk, rst, out_s3826, out_e3826, result3826);
PE P3827(out_s3763, out_e3826, clk, rst, out_s3827, out_e3827, result3827);
PE P3828(out_s3764, out_e3827, clk, rst, out_s3828, out_e3828, result3828);
PE P3829(out_s3765, out_e3828, clk, rst, out_s3829, out_e3829, result3829);
PE P3830(out_s3766, out_e3829, clk, rst, out_s3830, out_e3830, result3830);
PE P3831(out_s3767, out_e3830, clk, rst, out_s3831, out_e3831, result3831);
PE P3832(out_s3768, out_e3831, clk, rst, out_s3832, out_e3832, result3832);
PE P3833(out_s3769, out_e3832, clk, rst, out_s3833, out_e3833, result3833);
PE P3834(out_s3770, out_e3833, clk, rst, out_s3834, out_e3834, result3834);
PE P3835(out_s3771, out_e3834, clk, rst, out_s3835, out_e3835, result3835);
PE P3836(out_s3772, out_e3835, clk, rst, out_s3836, out_e3836, result3836);
PE P3837(out_s3773, out_e3836, clk, rst, out_s3837, out_e3837, result3837);
PE P3838(out_s3774, out_e3837, clk, rst, out_s3838, out_e3838, result3838);
PE P3839(out_s3775, out_e3838, clk, rst, out_s3839, out_e3839, result3839);

PE P3841(out_s3777, out_e3840, clk, rst, out_s3841, out_e3841, result3841);
PE P3842(out_s3778, out_e3841, clk, rst, out_s3842, out_e3842, result3842);
PE P3843(out_s3779, out_e3842, clk, rst, out_s3843, out_e3843, result3843);
PE P3844(out_s3780, out_e3843, clk, rst, out_s3844, out_e3844, result3844);
PE P3845(out_s3781, out_e3844, clk, rst, out_s3845, out_e3845, result3845);
PE P3846(out_s3782, out_e3845, clk, rst, out_s3846, out_e3846, result3846);
PE P3847(out_s3783, out_e3846, clk, rst, out_s3847, out_e3847, result3847);
PE P3848(out_s3784, out_e3847, clk, rst, out_s3848, out_e3848, result3848);
PE P3849(out_s3785, out_e3848, clk, rst, out_s3849, out_e3849, result3849);
PE P3850(out_s3786, out_e3849, clk, rst, out_s3850, out_e3850, result3850);
PE P3851(out_s3787, out_e3850, clk, rst, out_s3851, out_e3851, result3851);
PE P3852(out_s3788, out_e3851, clk, rst, out_s3852, out_e3852, result3852);
PE P3853(out_s3789, out_e3852, clk, rst, out_s3853, out_e3853, result3853);
PE P3854(out_s3790, out_e3853, clk, rst, out_s3854, out_e3854, result3854);
PE P3855(out_s3791, out_e3854, clk, rst, out_s3855, out_e3855, result3855);
PE P3856(out_s3792, out_e3855, clk, rst, out_s3856, out_e3856, result3856);
PE P3857(out_s3793, out_e3856, clk, rst, out_s3857, out_e3857, result3857);
PE P3858(out_s3794, out_e3857, clk, rst, out_s3858, out_e3858, result3858);
PE P3859(out_s3795, out_e3858, clk, rst, out_s3859, out_e3859, result3859);
PE P3860(out_s3796, out_e3859, clk, rst, out_s3860, out_e3860, result3860);
PE P3861(out_s3797, out_e3860, clk, rst, out_s3861, out_e3861, result3861);
PE P3862(out_s3798, out_e3861, clk, rst, out_s3862, out_e3862, result3862);
PE P3863(out_s3799, out_e3862, clk, rst, out_s3863, out_e3863, result3863);
PE P3864(out_s3800, out_e3863, clk, rst, out_s3864, out_e3864, result3864);
PE P3865(out_s3801, out_e3864, clk, rst, out_s3865, out_e3865, result3865);
PE P3866(out_s3802, out_e3865, clk, rst, out_s3866, out_e3866, result3866);
PE P3867(out_s3803, out_e3866, clk, rst, out_s3867, out_e3867, result3867);
PE P3868(out_s3804, out_e3867, clk, rst, out_s3868, out_e3868, result3868);
PE P3869(out_s3805, out_e3868, clk, rst, out_s3869, out_e3869, result3869);
PE P3870(out_s3806, out_e3869, clk, rst, out_s3870, out_e3870, result3870);
PE P3871(out_s3807, out_e3870, clk, rst, out_s3871, out_e3871, result3871);
PE P3872(out_s3808, out_e3871, clk, rst, out_s3872, out_e3872, result3872);
PE P3873(out_s3809, out_e3872, clk, rst, out_s3873, out_e3873, result3873);
PE P3874(out_s3810, out_e3873, clk, rst, out_s3874, out_e3874, result3874);
PE P3875(out_s3811, out_e3874, clk, rst, out_s3875, out_e3875, result3875);
PE P3876(out_s3812, out_e3875, clk, rst, out_s3876, out_e3876, result3876);
PE P3877(out_s3813, out_e3876, clk, rst, out_s3877, out_e3877, result3877);
PE P3878(out_s3814, out_e3877, clk, rst, out_s3878, out_e3878, result3878);
PE P3879(out_s3815, out_e3878, clk, rst, out_s3879, out_e3879, result3879);
PE P3880(out_s3816, out_e3879, clk, rst, out_s3880, out_e3880, result3880);
PE P3881(out_s3817, out_e3880, clk, rst, out_s3881, out_e3881, result3881);
PE P3882(out_s3818, out_e3881, clk, rst, out_s3882, out_e3882, result3882);
PE P3883(out_s3819, out_e3882, clk, rst, out_s3883, out_e3883, result3883);
PE P3884(out_s3820, out_e3883, clk, rst, out_s3884, out_e3884, result3884);
PE P3885(out_s3821, out_e3884, clk, rst, out_s3885, out_e3885, result3885);
PE P3886(out_s3822, out_e3885, clk, rst, out_s3886, out_e3886, result3886);
PE P3887(out_s3823, out_e3886, clk, rst, out_s3887, out_e3887, result3887);
PE P3888(out_s3824, out_e3887, clk, rst, out_s3888, out_e3888, result3888);
PE P3889(out_s3825, out_e3888, clk, rst, out_s3889, out_e3889, result3889);
PE P3890(out_s3826, out_e3889, clk, rst, out_s3890, out_e3890, result3890);
PE P3891(out_s3827, out_e3890, clk, rst, out_s3891, out_e3891, result3891);
PE P3892(out_s3828, out_e3891, clk, rst, out_s3892, out_e3892, result3892);
PE P3893(out_s3829, out_e3892, clk, rst, out_s3893, out_e3893, result3893);
PE P3894(out_s3830, out_e3893, clk, rst, out_s3894, out_e3894, result3894);
PE P3895(out_s3831, out_e3894, clk, rst, out_s3895, out_e3895, result3895);
PE P3896(out_s3832, out_e3895, clk, rst, out_s3896, out_e3896, result3896);
PE P3897(out_s3833, out_e3896, clk, rst, out_s3897, out_e3897, result3897);
PE P3898(out_s3834, out_e3897, clk, rst, out_s3898, out_e3898, result3898);
PE P3899(out_s3835, out_e3898, clk, rst, out_s3899, out_e3899, result3899);
PE P3900(out_s3836, out_e3899, clk, rst, out_s3900, out_e3900, result3900);
PE P3901(out_s3837, out_e3900, clk, rst, out_s3901, out_e3901, result3901);
PE P3902(out_s3838, out_e3901, clk, rst, out_s3902, out_e3902, result3902);
PE P3903(out_s3839, out_e3902, clk, rst, out_s3903, out_e3903, result3903);

PE P3905(out_s3841, out_e3904, clk, rst, out_s3905, out_e3905, result3905);
PE P3906(out_s3842, out_e3905, clk, rst, out_s3906, out_e3906, result3906);
PE P3907(out_s3843, out_e3906, clk, rst, out_s3907, out_e3907, result3907);
PE P3908(out_s3844, out_e3907, clk, rst, out_s3908, out_e3908, result3908);
PE P3909(out_s3845, out_e3908, clk, rst, out_s3909, out_e3909, result3909);
PE P3910(out_s3846, out_e3909, clk, rst, out_s3910, out_e3910, result3910);
PE P3911(out_s3847, out_e3910, clk, rst, out_s3911, out_e3911, result3911);
PE P3912(out_s3848, out_e3911, clk, rst, out_s3912, out_e3912, result3912);
PE P3913(out_s3849, out_e3912, clk, rst, out_s3913, out_e3913, result3913);
PE P3914(out_s3850, out_e3913, clk, rst, out_s3914, out_e3914, result3914);
PE P3915(out_s3851, out_e3914, clk, rst, out_s3915, out_e3915, result3915);
PE P3916(out_s3852, out_e3915, clk, rst, out_s3916, out_e3916, result3916);
PE P3917(out_s3853, out_e3916, clk, rst, out_s3917, out_e3917, result3917);
PE P3918(out_s3854, out_e3917, clk, rst, out_s3918, out_e3918, result3918);
PE P3919(out_s3855, out_e3918, clk, rst, out_s3919, out_e3919, result3919);
PE P3920(out_s3856, out_e3919, clk, rst, out_s3920, out_e3920, result3920);
PE P3921(out_s3857, out_e3920, clk, rst, out_s3921, out_e3921, result3921);
PE P3922(out_s3858, out_e3921, clk, rst, out_s3922, out_e3922, result3922);
PE P3923(out_s3859, out_e3922, clk, rst, out_s3923, out_e3923, result3923);
PE P3924(out_s3860, out_e3923, clk, rst, out_s3924, out_e3924, result3924);
PE P3925(out_s3861, out_e3924, clk, rst, out_s3925, out_e3925, result3925);
PE P3926(out_s3862, out_e3925, clk, rst, out_s3926, out_e3926, result3926);
PE P3927(out_s3863, out_e3926, clk, rst, out_s3927, out_e3927, result3927);
PE P3928(out_s3864, out_e3927, clk, rst, out_s3928, out_e3928, result3928);
PE P3929(out_s3865, out_e3928, clk, rst, out_s3929, out_e3929, result3929);
PE P3930(out_s3866, out_e3929, clk, rst, out_s3930, out_e3930, result3930);
PE P3931(out_s3867, out_e3930, clk, rst, out_s3931, out_e3931, result3931);
PE P3932(out_s3868, out_e3931, clk, rst, out_s3932, out_e3932, result3932);
PE P3933(out_s3869, out_e3932, clk, rst, out_s3933, out_e3933, result3933);
PE P3934(out_s3870, out_e3933, clk, rst, out_s3934, out_e3934, result3934);
PE P3935(out_s3871, out_e3934, clk, rst, out_s3935, out_e3935, result3935);
PE P3936(out_s3872, out_e3935, clk, rst, out_s3936, out_e3936, result3936);
PE P3937(out_s3873, out_e3936, clk, rst, out_s3937, out_e3937, result3937);
PE P3938(out_s3874, out_e3937, clk, rst, out_s3938, out_e3938, result3938);
PE P3939(out_s3875, out_e3938, clk, rst, out_s3939, out_e3939, result3939);
PE P3940(out_s3876, out_e3939, clk, rst, out_s3940, out_e3940, result3940);
PE P3941(out_s3877, out_e3940, clk, rst, out_s3941, out_e3941, result3941);
PE P3942(out_s3878, out_e3941, clk, rst, out_s3942, out_e3942, result3942);
PE P3943(out_s3879, out_e3942, clk, rst, out_s3943, out_e3943, result3943);
PE P3944(out_s3880, out_e3943, clk, rst, out_s3944, out_e3944, result3944);
PE P3945(out_s3881, out_e3944, clk, rst, out_s3945, out_e3945, result3945);
PE P3946(out_s3882, out_e3945, clk, rst, out_s3946, out_e3946, result3946);
PE P3947(out_s3883, out_e3946, clk, rst, out_s3947, out_e3947, result3947);
PE P3948(out_s3884, out_e3947, clk, rst, out_s3948, out_e3948, result3948);
PE P3949(out_s3885, out_e3948, clk, rst, out_s3949, out_e3949, result3949);
PE P3950(out_s3886, out_e3949, clk, rst, out_s3950, out_e3950, result3950);
PE P3951(out_s3887, out_e3950, clk, rst, out_s3951, out_e3951, result3951);
PE P3952(out_s3888, out_e3951, clk, rst, out_s3952, out_e3952, result3952);
PE P3953(out_s3889, out_e3952, clk, rst, out_s3953, out_e3953, result3953);
PE P3954(out_s3890, out_e3953, clk, rst, out_s3954, out_e3954, result3954);
PE P3955(out_s3891, out_e3954, clk, rst, out_s3955, out_e3955, result3955);
PE P3956(out_s3892, out_e3955, clk, rst, out_s3956, out_e3956, result3956);
PE P3957(out_s3893, out_e3956, clk, rst, out_s3957, out_e3957, result3957);
PE P3958(out_s3894, out_e3957, clk, rst, out_s3958, out_e3958, result3958);
PE P3959(out_s3895, out_e3958, clk, rst, out_s3959, out_e3959, result3959);
PE P3960(out_s3896, out_e3959, clk, rst, out_s3960, out_e3960, result3960);
PE P3961(out_s3897, out_e3960, clk, rst, out_s3961, out_e3961, result3961);
PE P3962(out_s3898, out_e3961, clk, rst, out_s3962, out_e3962, result3962);
PE P3963(out_s3899, out_e3962, clk, rst, out_s3963, out_e3963, result3963);
PE P3964(out_s3900, out_e3963, clk, rst, out_s3964, out_e3964, result3964);
PE P3965(out_s3901, out_e3964, clk, rst, out_s3965, out_e3965, result3965);
PE P3966(out_s3902, out_e3965, clk, rst, out_s3966, out_e3966, result3966);
PE P3967(out_s3903, out_e3966, clk, rst, out_s3967, out_e3967, result3967);

PE P3969(out_s3905, out_e3968, clk, rst, out_s3969, out_e3969, result3969);
PE P3970(out_s3906, out_e3969, clk, rst, out_s3970, out_e3970, result3970);
PE P3971(out_s3907, out_e3970, clk, rst, out_s3971, out_e3971, result3971);
PE P3972(out_s3908, out_e3971, clk, rst, out_s3972, out_e3972, result3972);
PE P3973(out_s3909, out_e3972, clk, rst, out_s3973, out_e3973, result3973);
PE P3974(out_s3910, out_e3973, clk, rst, out_s3974, out_e3974, result3974);
PE P3975(out_s3911, out_e3974, clk, rst, out_s3975, out_e3975, result3975);
PE P3976(out_s3912, out_e3975, clk, rst, out_s3976, out_e3976, result3976);
PE P3977(out_s3913, out_e3976, clk, rst, out_s3977, out_e3977, result3977);
PE P3978(out_s3914, out_e3977, clk, rst, out_s3978, out_e3978, result3978);
PE P3979(out_s3915, out_e3978, clk, rst, out_s3979, out_e3979, result3979);
PE P3980(out_s3916, out_e3979, clk, rst, out_s3980, out_e3980, result3980);
PE P3981(out_s3917, out_e3980, clk, rst, out_s3981, out_e3981, result3981);
PE P3982(out_s3918, out_e3981, clk, rst, out_s3982, out_e3982, result3982);
PE P3983(out_s3919, out_e3982, clk, rst, out_s3983, out_e3983, result3983);
PE P3984(out_s3920, out_e3983, clk, rst, out_s3984, out_e3984, result3984);
PE P3985(out_s3921, out_e3984, clk, rst, out_s3985, out_e3985, result3985);
PE P3986(out_s3922, out_e3985, clk, rst, out_s3986, out_e3986, result3986);
PE P3987(out_s3923, out_e3986, clk, rst, out_s3987, out_e3987, result3987);
PE P3988(out_s3924, out_e3987, clk, rst, out_s3988, out_e3988, result3988);
PE P3989(out_s3925, out_e3988, clk, rst, out_s3989, out_e3989, result3989);
PE P3990(out_s3926, out_e3989, clk, rst, out_s3990, out_e3990, result3990);
PE P3991(out_s3927, out_e3990, clk, rst, out_s3991, out_e3991, result3991);
PE P3992(out_s3928, out_e3991, clk, rst, out_s3992, out_e3992, result3992);
PE P3993(out_s3929, out_e3992, clk, rst, out_s3993, out_e3993, result3993);
PE P3994(out_s3930, out_e3993, clk, rst, out_s3994, out_e3994, result3994);
PE P3995(out_s3931, out_e3994, clk, rst, out_s3995, out_e3995, result3995);
PE P3996(out_s3932, out_e3995, clk, rst, out_s3996, out_e3996, result3996);
PE P3997(out_s3933, out_e3996, clk, rst, out_s3997, out_e3997, result3997);
PE P3998(out_s3934, out_e3997, clk, rst, out_s3998, out_e3998, result3998);
PE P3999(out_s3935, out_e3998, clk, rst, out_s3999, out_e3999, result3999);
PE P4000(out_s3936, out_e3999, clk, rst, out_s4000, out_e4000, result4000);
PE P4001(out_s3937, out_e4000, clk, rst, out_s4001, out_e4001, result4001);
PE P4002(out_s3938, out_e4001, clk, rst, out_s4002, out_e4002, result4002);
PE P4003(out_s3939, out_e4002, clk, rst, out_s4003, out_e4003, result4003);
PE P4004(out_s3940, out_e4003, clk, rst, out_s4004, out_e4004, result4004);
PE P4005(out_s3941, out_e4004, clk, rst, out_s4005, out_e4005, result4005);
PE P4006(out_s3942, out_e4005, clk, rst, out_s4006, out_e4006, result4006);
PE P4007(out_s3943, out_e4006, clk, rst, out_s4007, out_e4007, result4007);
PE P4008(out_s3944, out_e4007, clk, rst, out_s4008, out_e4008, result4008);
PE P4009(out_s3945, out_e4008, clk, rst, out_s4009, out_e4009, result4009);
PE P4010(out_s3946, out_e4009, clk, rst, out_s4010, out_e4010, result4010);
PE P4011(out_s3947, out_e4010, clk, rst, out_s4011, out_e4011, result4011);
PE P4012(out_s3948, out_e4011, clk, rst, out_s4012, out_e4012, result4012);
PE P4013(out_s3949, out_e4012, clk, rst, out_s4013, out_e4013, result4013);
PE P4014(out_s3950, out_e4013, clk, rst, out_s4014, out_e4014, result4014);
PE P4015(out_s3951, out_e4014, clk, rst, out_s4015, out_e4015, result4015);
PE P4016(out_s3952, out_e4015, clk, rst, out_s4016, out_e4016, result4016);
PE P4017(out_s3953, out_e4016, clk, rst, out_s4017, out_e4017, result4017);
PE P4018(out_s3954, out_e4017, clk, rst, out_s4018, out_e4018, result4018);
PE P4019(out_s3955, out_e4018, clk, rst, out_s4019, out_e4019, result4019);
PE P4020(out_s3956, out_e4019, clk, rst, out_s4020, out_e4020, result4020);
PE P4021(out_s3957, out_e4020, clk, rst, out_s4021, out_e4021, result4021);
PE P4022(out_s3958, out_e4021, clk, rst, out_s4022, out_e4022, result4022);
PE P4023(out_s3959, out_e4022, clk, rst, out_s4023, out_e4023, result4023);
PE P4024(out_s3960, out_e4023, clk, rst, out_s4024, out_e4024, result4024);
PE P4025(out_s3961, out_e4024, clk, rst, out_s4025, out_e4025, result4025);
PE P4026(out_s3962, out_e4025, clk, rst, out_s4026, out_e4026, result4026);
PE P4027(out_s3963, out_e4026, clk, rst, out_s4027, out_e4027, result4027);
PE P4028(out_s3964, out_e4027, clk, rst, out_s4028, out_e4028, result4028);
PE P4029(out_s3965, out_e4028, clk, rst, out_s4029, out_e4029, result4029);
PE P4030(out_s3966, out_e4029, clk, rst, out_s4030, out_e4030, result4030);
PE P4031(out_s3967, out_e4030, clk, rst, out_s4031, out_e4031, result4031);

PE P4033(out_s3969, out_e4032, clk, rst, out_s4033, out_e4033, result4033);
PE P4034(out_s3970, out_e4033, clk, rst, out_s4034, out_e4034, result4034);
PE P4035(out_s3971, out_e4034, clk, rst, out_s4035, out_e4035, result4035);
PE P4036(out_s3972, out_e4035, clk, rst, out_s4036, out_e4036, result4036);
PE P4037(out_s3973, out_e4036, clk, rst, out_s4037, out_e4037, result4037);
PE P4038(out_s3974, out_e4037, clk, rst, out_s4038, out_e4038, result4038);
PE P4039(out_s3975, out_e4038, clk, rst, out_s4039, out_e4039, result4039);
PE P4040(out_s3976, out_e4039, clk, rst, out_s4040, out_e4040, result4040);
PE P4041(out_s3977, out_e4040, clk, rst, out_s4041, out_e4041, result4041);
PE P4042(out_s3978, out_e4041, clk, rst, out_s4042, out_e4042, result4042);
PE P4043(out_s3979, out_e4042, clk, rst, out_s4043, out_e4043, result4043);
PE P4044(out_s3980, out_e4043, clk, rst, out_s4044, out_e4044, result4044);
PE P4045(out_s3981, out_e4044, clk, rst, out_s4045, out_e4045, result4045);
PE P4046(out_s3982, out_e4045, clk, rst, out_s4046, out_e4046, result4046);
PE P4047(out_s3983, out_e4046, clk, rst, out_s4047, out_e4047, result4047);
PE P4048(out_s3984, out_e4047, clk, rst, out_s4048, out_e4048, result4048);
PE P4049(out_s3985, out_e4048, clk, rst, out_s4049, out_e4049, result4049);
PE P4050(out_s3986, out_e4049, clk, rst, out_s4050, out_e4050, result4050);
PE P4051(out_s3987, out_e4050, clk, rst, out_s4051, out_e4051, result4051);
PE P4052(out_s3988, out_e4051, clk, rst, out_s4052, out_e4052, result4052);
PE P4053(out_s3989, out_e4052, clk, rst, out_s4053, out_e4053, result4053);
PE P4054(out_s3990, out_e4053, clk, rst, out_s4054, out_e4054, result4054);
PE P4055(out_s3991, out_e4054, clk, rst, out_s4055, out_e4055, result4055);
PE P4056(out_s3992, out_e4055, clk, rst, out_s4056, out_e4056, result4056);
PE P4057(out_s3993, out_e4056, clk, rst, out_s4057, out_e4057, result4057);
PE P4058(out_s3994, out_e4057, clk, rst, out_s4058, out_e4058, result4058);
PE P4059(out_s3995, out_e4058, clk, rst, out_s4059, out_e4059, result4059);
PE P4060(out_s3996, out_e4059, clk, rst, out_s4060, out_e4060, result4060);
PE P4061(out_s3997, out_e4060, clk, rst, out_s4061, out_e4061, result4061);
PE P4062(out_s3998, out_e4061, clk, rst, out_s4062, out_e4062, result4062);
PE P4063(out_s3999, out_e4062, clk, rst, out_s4063, out_e4063, result4063);
PE P4064(out_s4000, out_e4063, clk, rst, out_s4064, out_e4064, result4064);
PE P4065(out_s4001, out_e4064, clk, rst, out_s4065, out_e4065, result4065);
PE P4066(out_s4002, out_e4065, clk, rst, out_s4066, out_e4066, result4066);
PE P4067(out_s4003, out_e4066, clk, rst, out_s4067, out_e4067, result4067);
PE P4068(out_s4004, out_e4067, clk, rst, out_s4068, out_e4068, result4068);
PE P4069(out_s4005, out_e4068, clk, rst, out_s4069, out_e4069, result4069);
PE P4070(out_s4006, out_e4069, clk, rst, out_s4070, out_e4070, result4070);
PE P4071(out_s4007, out_e4070, clk, rst, out_s4071, out_e4071, result4071);
PE P4072(out_s4008, out_e4071, clk, rst, out_s4072, out_e4072, result4072);
PE P4073(out_s4009, out_e4072, clk, rst, out_s4073, out_e4073, result4073);
PE P4074(out_s4010, out_e4073, clk, rst, out_s4074, out_e4074, result4074);
PE P4075(out_s4011, out_e4074, clk, rst, out_s4075, out_e4075, result4075);
PE P4076(out_s4012, out_e4075, clk, rst, out_s4076, out_e4076, result4076);
PE P4077(out_s4013, out_e4076, clk, rst, out_s4077, out_e4077, result4077);
PE P4078(out_s4014, out_e4077, clk, rst, out_s4078, out_e4078, result4078);
PE P4079(out_s4015, out_e4078, clk, rst, out_s4079, out_e4079, result4079);
PE P4080(out_s4016, out_e4079, clk, rst, out_s4080, out_e4080, result4080);
PE P4081(out_s4017, out_e4080, clk, rst, out_s4081, out_e4081, result4081);
PE P4082(out_s4018, out_e4081, clk, rst, out_s4082, out_e4082, result4082);
PE P4083(out_s4019, out_e4082, clk, rst, out_s4083, out_e4083, result4083);
PE P4084(out_s4020, out_e4083, clk, rst, out_s4084, out_e4084, result4084);
PE P4085(out_s4021, out_e4084, clk, rst, out_s4085, out_e4085, result4085);
PE P4086(out_s4022, out_e4085, clk, rst, out_s4086, out_e4086, result4086);
PE P4087(out_s4023, out_e4086, clk, rst, out_s4087, out_e4087, result4087);
PE P4088(out_s4024, out_e4087, clk, rst, out_s4088, out_e4088, result4088);
PE P4089(out_s4025, out_e4088, clk, rst, out_s4089, out_e4089, result4089);
PE P4090(out_s4026, out_e4089, clk, rst, out_s4090, out_e4090, result4090);
PE P4091(out_s4027, out_e4090, clk, rst, out_s4091, out_e4091, result4091);
PE P4092(out_s4028, out_e4091, clk, rst, out_s4092, out_e4092, result4092);
PE P4093(out_s4029, out_e4092, clk, rst, out_s4093, out_e4093, result4093);
PE P4094(out_s4030, out_e4093, clk, rst, out_s4094, out_e4094, result4094);
PE P4095(out_s4031, out_e4094, clk, rst, out_s4095, out_e4095, result4095);

always @(posedge clk or posedge rst) begin
    if(rst) begin
        done <= 0;
        count <= 0;
    end
    else begin
		result_out0<=result0;
		result_out1<=result1;
		result_out2<=result2;
		result_out3<=result3;
		result_out4<=result4;
		result_out5<=result5;
		result_out6<=result6;
		result_out7<=result7;
		result_out8<=result8;
		result_out9<=result9;
		result_out10<=result10;
		result_out11<=result11;
		result_out12<=result12;
		result_out13<=result13;
		result_out14<=result14;
		result_out15<=result15;
		result_out16<=result16;
		result_out17<=result17;
		result_out18<=result18;
		result_out19<=result19;
		result_out20<=result20;
		result_out21<=result21;
		result_out22<=result22;
		result_out23<=result23;
		result_out24<=result24;
		result_out25<=result25;
		result_out26<=result26;
		result_out27<=result27;
		result_out28<=result28;
		result_out29<=result29;
		result_out30<=result30;
		result_out31<=result31;
		result_out32<=result32;
		result_out33<=result33;
		result_out34<=result34;
		result_out35<=result35;
		result_out36<=result36;
		result_out37<=result37;
		result_out38<=result38;
		result_out39<=result39;
		result_out40<=result40;
		result_out41<=result41;
		result_out42<=result42;
		result_out43<=result43;
		result_out44<=result44;
		result_out45<=result45;
		result_out46<=result46;
		result_out47<=result47;
		result_out48<=result48;
		result_out49<=result49;
		result_out50<=result50;
		result_out51<=result51;
		result_out52<=result52;
		result_out53<=result53;
		result_out54<=result54;
		result_out55<=result55;
		result_out56<=result56;
		result_out57<=result57;
		result_out58<=result58;
		result_out59<=result59;
		result_out60<=result60;
		result_out61<=result61;
		result_out62<=result62;
		result_out63<=result63;
		result_out64<=result64;
		result_out65<=result65;
		result_out66<=result66;
		result_out67<=result67;
		result_out68<=result68;
		result_out69<=result69;
		result_out70<=result70;
		result_out71<=result71;
		result_out72<=result72;
		result_out73<=result73;
		result_out74<=result74;
		result_out75<=result75;
		result_out76<=result76;
		result_out77<=result77;
		result_out78<=result78;
		result_out79<=result79;
		result_out80<=result80;
		result_out81<=result81;
		result_out82<=result82;
		result_out83<=result83;
		result_out84<=result84;
		result_out85<=result85;
		result_out86<=result86;
		result_out87<=result87;
		result_out88<=result88;
		result_out89<=result89;
		result_out90<=result90;
		result_out91<=result91;
		result_out92<=result92;
		result_out93<=result93;
		result_out94<=result94;
		result_out95<=result95;
		result_out96<=result96;
		result_out97<=result97;
		result_out98<=result98;
		result_out99<=result99;
		result_out100<=result100;
		result_out101<=result101;
		result_out102<=result102;
		result_out103<=result103;
		result_out104<=result104;
		result_out105<=result105;
		result_out106<=result106;
		result_out107<=result107;
		result_out108<=result108;
		result_out109<=result109;
		result_out110<=result110;
		result_out111<=result111;
		result_out112<=result112;
		result_out113<=result113;
		result_out114<=result114;
		result_out115<=result115;
		result_out116<=result116;
		result_out117<=result117;
		result_out118<=result118;
		result_out119<=result119;
		result_out120<=result120;
		result_out121<=result121;
		result_out122<=result122;
		result_out123<=result123;
		result_out124<=result124;
		result_out125<=result125;
		result_out126<=result126;
		result_out127<=result127;
		result_out128<=result128;
		result_out129<=result129;
		result_out130<=result130;
		result_out131<=result131;
		result_out132<=result132;
		result_out133<=result133;
		result_out134<=result134;
		result_out135<=result135;
		result_out136<=result136;
		result_out137<=result137;
		result_out138<=result138;
		result_out139<=result139;
		result_out140<=result140;
		result_out141<=result141;
		result_out142<=result142;
		result_out143<=result143;
		result_out144<=result144;
		result_out145<=result145;
		result_out146<=result146;
		result_out147<=result147;
		result_out148<=result148;
		result_out149<=result149;
		result_out150<=result150;
		result_out151<=result151;
		result_out152<=result152;
		result_out153<=result153;
		result_out154<=result154;
		result_out155<=result155;
		result_out156<=result156;
		result_out157<=result157;
		result_out158<=result158;
		result_out159<=result159;
		result_out160<=result160;
		result_out161<=result161;
		result_out162<=result162;
		result_out163<=result163;
		result_out164<=result164;
		result_out165<=result165;
		result_out166<=result166;
		result_out167<=result167;
		result_out168<=result168;
		result_out169<=result169;
		result_out170<=result170;
		result_out171<=result171;
		result_out172<=result172;
		result_out173<=result173;
		result_out174<=result174;
		result_out175<=result175;
		result_out176<=result176;
		result_out177<=result177;
		result_out178<=result178;
		result_out179<=result179;
		result_out180<=result180;
		result_out181<=result181;
		result_out182<=result182;
		result_out183<=result183;
		result_out184<=result184;
		result_out185<=result185;
		result_out186<=result186;
		result_out187<=result187;
		result_out188<=result188;
		result_out189<=result189;
		result_out190<=result190;
		result_out191<=result191;
		result_out192<=result192;
		result_out193<=result193;
		result_out194<=result194;
		result_out195<=result195;
		result_out196<=result196;
		result_out197<=result197;
		result_out198<=result198;
		result_out199<=result199;
		result_out200<=result200;
		result_out201<=result201;
		result_out202<=result202;
		result_out203<=result203;
		result_out204<=result204;
		result_out205<=result205;
		result_out206<=result206;
		result_out207<=result207;
		result_out208<=result208;
		result_out209<=result209;
		result_out210<=result210;
		result_out211<=result211;
		result_out212<=result212;
		result_out213<=result213;
		result_out214<=result214;
		result_out215<=result215;
		result_out216<=result216;
		result_out217<=result217;
		result_out218<=result218;
		result_out219<=result219;
		result_out220<=result220;
		result_out221<=result221;
		result_out222<=result222;
		result_out223<=result223;
		result_out224<=result224;
		result_out225<=result225;
		result_out226<=result226;
		result_out227<=result227;
		result_out228<=result228;
		result_out229<=result229;
		result_out230<=result230;
		result_out231<=result231;
		result_out232<=result232;
		result_out233<=result233;
		result_out234<=result234;
		result_out235<=result235;
		result_out236<=result236;
		result_out237<=result237;
		result_out238<=result238;
		result_out239<=result239;
		result_out240<=result240;
		result_out241<=result241;
		result_out242<=result242;
		result_out243<=result243;
		result_out244<=result244;
		result_out245<=result245;
		result_out246<=result246;
		result_out247<=result247;
		result_out248<=result248;
		result_out249<=result249;
		result_out250<=result250;
		result_out251<=result251;
		result_out252<=result252;
		result_out253<=result253;
		result_out254<=result254;
		result_out255<=result255;
		result_out256<=result256;
		result_out257<=result257;
		result_out258<=result258;
		result_out259<=result259;
		result_out260<=result260;
		result_out261<=result261;
		result_out262<=result262;
		result_out263<=result263;
		result_out264<=result264;
		result_out265<=result265;
		result_out266<=result266;
		result_out267<=result267;
		result_out268<=result268;
		result_out269<=result269;
		result_out270<=result270;
		result_out271<=result271;
		result_out272<=result272;
		result_out273<=result273;
		result_out274<=result274;
		result_out275<=result275;
		result_out276<=result276;
		result_out277<=result277;
		result_out278<=result278;
		result_out279<=result279;
		result_out280<=result280;
		result_out281<=result281;
		result_out282<=result282;
		result_out283<=result283;
		result_out284<=result284;
		result_out285<=result285;
		result_out286<=result286;
		result_out287<=result287;
		result_out288<=result288;
		result_out289<=result289;
		result_out290<=result290;
		result_out291<=result291;
		result_out292<=result292;
		result_out293<=result293;
		result_out294<=result294;
		result_out295<=result295;
		result_out296<=result296;
		result_out297<=result297;
		result_out298<=result298;
		result_out299<=result299;
		result_out300<=result300;
		result_out301<=result301;
		result_out302<=result302;
		result_out303<=result303;
		result_out304<=result304;
		result_out305<=result305;
		result_out306<=result306;
		result_out307<=result307;
		result_out308<=result308;
		result_out309<=result309;
		result_out310<=result310;
		result_out311<=result311;
		result_out312<=result312;
		result_out313<=result313;
		result_out314<=result314;
		result_out315<=result315;
		result_out316<=result316;
		result_out317<=result317;
		result_out318<=result318;
		result_out319<=result319;
		result_out320<=result320;
		result_out321<=result321;
		result_out322<=result322;
		result_out323<=result323;
		result_out324<=result324;
		result_out325<=result325;
		result_out326<=result326;
		result_out327<=result327;
		result_out328<=result328;
		result_out329<=result329;
		result_out330<=result330;
		result_out331<=result331;
		result_out332<=result332;
		result_out333<=result333;
		result_out334<=result334;
		result_out335<=result335;
		result_out336<=result336;
		result_out337<=result337;
		result_out338<=result338;
		result_out339<=result339;
		result_out340<=result340;
		result_out341<=result341;
		result_out342<=result342;
		result_out343<=result343;
		result_out344<=result344;
		result_out345<=result345;
		result_out346<=result346;
		result_out347<=result347;
		result_out348<=result348;
		result_out349<=result349;
		result_out350<=result350;
		result_out351<=result351;
		result_out352<=result352;
		result_out353<=result353;
		result_out354<=result354;
		result_out355<=result355;
		result_out356<=result356;
		result_out357<=result357;
		result_out358<=result358;
		result_out359<=result359;
		result_out360<=result360;
		result_out361<=result361;
		result_out362<=result362;
		result_out363<=result363;
		result_out364<=result364;
		result_out365<=result365;
		result_out366<=result366;
		result_out367<=result367;
		result_out368<=result368;
		result_out369<=result369;
		result_out370<=result370;
		result_out371<=result371;
		result_out372<=result372;
		result_out373<=result373;
		result_out374<=result374;
		result_out375<=result375;
		result_out376<=result376;
		result_out377<=result377;
		result_out378<=result378;
		result_out379<=result379;
		result_out380<=result380;
		result_out381<=result381;
		result_out382<=result382;
		result_out383<=result383;
		result_out384<=result384;
		result_out385<=result385;
		result_out386<=result386;
		result_out387<=result387;
		result_out388<=result388;
		result_out389<=result389;
		result_out390<=result390;
		result_out391<=result391;
		result_out392<=result392;
		result_out393<=result393;
		result_out394<=result394;
		result_out395<=result395;
		result_out396<=result396;
		result_out397<=result397;
		result_out398<=result398;
		result_out399<=result399;
		result_out400<=result400;
		result_out401<=result401;
		result_out402<=result402;
		result_out403<=result403;
		result_out404<=result404;
		result_out405<=result405;
		result_out406<=result406;
		result_out407<=result407;
		result_out408<=result408;
		result_out409<=result409;
		result_out410<=result410;
		result_out411<=result411;
		result_out412<=result412;
		result_out413<=result413;
		result_out414<=result414;
		result_out415<=result415;
		result_out416<=result416;
		result_out417<=result417;
		result_out418<=result418;
		result_out419<=result419;
		result_out420<=result420;
		result_out421<=result421;
		result_out422<=result422;
		result_out423<=result423;
		result_out424<=result424;
		result_out425<=result425;
		result_out426<=result426;
		result_out427<=result427;
		result_out428<=result428;
		result_out429<=result429;
		result_out430<=result430;
		result_out431<=result431;
		result_out432<=result432;
		result_out433<=result433;
		result_out434<=result434;
		result_out435<=result435;
		result_out436<=result436;
		result_out437<=result437;
		result_out438<=result438;
		result_out439<=result439;
		result_out440<=result440;
		result_out441<=result441;
		result_out442<=result442;
		result_out443<=result443;
		result_out444<=result444;
		result_out445<=result445;
		result_out446<=result446;
		result_out447<=result447;
		result_out448<=result448;
		result_out449<=result449;
		result_out450<=result450;
		result_out451<=result451;
		result_out452<=result452;
		result_out453<=result453;
		result_out454<=result454;
		result_out455<=result455;
		result_out456<=result456;
		result_out457<=result457;
		result_out458<=result458;
		result_out459<=result459;
		result_out460<=result460;
		result_out461<=result461;
		result_out462<=result462;
		result_out463<=result463;
		result_out464<=result464;
		result_out465<=result465;
		result_out466<=result466;
		result_out467<=result467;
		result_out468<=result468;
		result_out469<=result469;
		result_out470<=result470;
		result_out471<=result471;
		result_out472<=result472;
		result_out473<=result473;
		result_out474<=result474;
		result_out475<=result475;
		result_out476<=result476;
		result_out477<=result477;
		result_out478<=result478;
		result_out479<=result479;
		result_out480<=result480;
		result_out481<=result481;
		result_out482<=result482;
		result_out483<=result483;
		result_out484<=result484;
		result_out485<=result485;
		result_out486<=result486;
		result_out487<=result487;
		result_out488<=result488;
		result_out489<=result489;
		result_out490<=result490;
		result_out491<=result491;
		result_out492<=result492;
		result_out493<=result493;
		result_out494<=result494;
		result_out495<=result495;
		result_out496<=result496;
		result_out497<=result497;
		result_out498<=result498;
		result_out499<=result499;
		result_out500<=result500;
		result_out501<=result501;
		result_out502<=result502;
		result_out503<=result503;
		result_out504<=result504;
		result_out505<=result505;
		result_out506<=result506;
		result_out507<=result507;
		result_out508<=result508;
		result_out509<=result509;
		result_out510<=result510;
		result_out511<=result511;
		result_out512<=result512;
		result_out513<=result513;
		result_out514<=result514;
		result_out515<=result515;
		result_out516<=result516;
		result_out517<=result517;
		result_out518<=result518;
		result_out519<=result519;
		result_out520<=result520;
		result_out521<=result521;
		result_out522<=result522;
		result_out523<=result523;
		result_out524<=result524;
		result_out525<=result525;
		result_out526<=result526;
		result_out527<=result527;
		result_out528<=result528;
		result_out529<=result529;
		result_out530<=result530;
		result_out531<=result531;
		result_out532<=result532;
		result_out533<=result533;
		result_out534<=result534;
		result_out535<=result535;
		result_out536<=result536;
		result_out537<=result537;
		result_out538<=result538;
		result_out539<=result539;
		result_out540<=result540;
		result_out541<=result541;
		result_out542<=result542;
		result_out543<=result543;
		result_out544<=result544;
		result_out545<=result545;
		result_out546<=result546;
		result_out547<=result547;
		result_out548<=result548;
		result_out549<=result549;
		result_out550<=result550;
		result_out551<=result551;
		result_out552<=result552;
		result_out553<=result553;
		result_out554<=result554;
		result_out555<=result555;
		result_out556<=result556;
		result_out557<=result557;
		result_out558<=result558;
		result_out559<=result559;
		result_out560<=result560;
		result_out561<=result561;
		result_out562<=result562;
		result_out563<=result563;
		result_out564<=result564;
		result_out565<=result565;
		result_out566<=result566;
		result_out567<=result567;
		result_out568<=result568;
		result_out569<=result569;
		result_out570<=result570;
		result_out571<=result571;
		result_out572<=result572;
		result_out573<=result573;
		result_out574<=result574;
		result_out575<=result575;
		result_out576<=result576;
		result_out577<=result577;
		result_out578<=result578;
		result_out579<=result579;
		result_out580<=result580;
		result_out581<=result581;
		result_out582<=result582;
		result_out583<=result583;
		result_out584<=result584;
		result_out585<=result585;
		result_out586<=result586;
		result_out587<=result587;
		result_out588<=result588;
		result_out589<=result589;
		result_out590<=result590;
		result_out591<=result591;
		result_out592<=result592;
		result_out593<=result593;
		result_out594<=result594;
		result_out595<=result595;
		result_out596<=result596;
		result_out597<=result597;
		result_out598<=result598;
		result_out599<=result599;
		result_out600<=result600;
		result_out601<=result601;
		result_out602<=result602;
		result_out603<=result603;
		result_out604<=result604;
		result_out605<=result605;
		result_out606<=result606;
		result_out607<=result607;
		result_out608<=result608;
		result_out609<=result609;
		result_out610<=result610;
		result_out611<=result611;
		result_out612<=result612;
		result_out613<=result613;
		result_out614<=result614;
		result_out615<=result615;
		result_out616<=result616;
		result_out617<=result617;
		result_out618<=result618;
		result_out619<=result619;
		result_out620<=result620;
		result_out621<=result621;
		result_out622<=result622;
		result_out623<=result623;
		result_out624<=result624;
		result_out625<=result625;
		result_out626<=result626;
		result_out627<=result627;
		result_out628<=result628;
		result_out629<=result629;
		result_out630<=result630;
		result_out631<=result631;
		result_out632<=result632;
		result_out633<=result633;
		result_out634<=result634;
		result_out635<=result635;
		result_out636<=result636;
		result_out637<=result637;
		result_out638<=result638;
		result_out639<=result639;
		result_out640<=result640;
		result_out641<=result641;
		result_out642<=result642;
		result_out643<=result643;
		result_out644<=result644;
		result_out645<=result645;
		result_out646<=result646;
		result_out647<=result647;
		result_out648<=result648;
		result_out649<=result649;
		result_out650<=result650;
		result_out651<=result651;
		result_out652<=result652;
		result_out653<=result653;
		result_out654<=result654;
		result_out655<=result655;
		result_out656<=result656;
		result_out657<=result657;
		result_out658<=result658;
		result_out659<=result659;
		result_out660<=result660;
		result_out661<=result661;
		result_out662<=result662;
		result_out663<=result663;
		result_out664<=result664;
		result_out665<=result665;
		result_out666<=result666;
		result_out667<=result667;
		result_out668<=result668;
		result_out669<=result669;
		result_out670<=result670;
		result_out671<=result671;
		result_out672<=result672;
		result_out673<=result673;
		result_out674<=result674;
		result_out675<=result675;
		result_out676<=result676;
		result_out677<=result677;
		result_out678<=result678;
		result_out679<=result679;
		result_out680<=result680;
		result_out681<=result681;
		result_out682<=result682;
		result_out683<=result683;
		result_out684<=result684;
		result_out685<=result685;
		result_out686<=result686;
		result_out687<=result687;
		result_out688<=result688;
		result_out689<=result689;
		result_out690<=result690;
		result_out691<=result691;
		result_out692<=result692;
		result_out693<=result693;
		result_out694<=result694;
		result_out695<=result695;
		result_out696<=result696;
		result_out697<=result697;
		result_out698<=result698;
		result_out699<=result699;
		result_out700<=result700;
		result_out701<=result701;
		result_out702<=result702;
		result_out703<=result703;
		result_out704<=result704;
		result_out705<=result705;
		result_out706<=result706;
		result_out707<=result707;
		result_out708<=result708;
		result_out709<=result709;
		result_out710<=result710;
		result_out711<=result711;
		result_out712<=result712;
		result_out713<=result713;
		result_out714<=result714;
		result_out715<=result715;
		result_out716<=result716;
		result_out717<=result717;
		result_out718<=result718;
		result_out719<=result719;
		result_out720<=result720;
		result_out721<=result721;
		result_out722<=result722;
		result_out723<=result723;
		result_out724<=result724;
		result_out725<=result725;
		result_out726<=result726;
		result_out727<=result727;
		result_out728<=result728;
		result_out729<=result729;
		result_out730<=result730;
		result_out731<=result731;
		result_out732<=result732;
		result_out733<=result733;
		result_out734<=result734;
		result_out735<=result735;
		result_out736<=result736;
		result_out737<=result737;
		result_out738<=result738;
		result_out739<=result739;
		result_out740<=result740;
		result_out741<=result741;
		result_out742<=result742;
		result_out743<=result743;
		result_out744<=result744;
		result_out745<=result745;
		result_out746<=result746;
		result_out747<=result747;
		result_out748<=result748;
		result_out749<=result749;
		result_out750<=result750;
		result_out751<=result751;
		result_out752<=result752;
		result_out753<=result753;
		result_out754<=result754;
		result_out755<=result755;
		result_out756<=result756;
		result_out757<=result757;
		result_out758<=result758;
		result_out759<=result759;
		result_out760<=result760;
		result_out761<=result761;
		result_out762<=result762;
		result_out763<=result763;
		result_out764<=result764;
		result_out765<=result765;
		result_out766<=result766;
		result_out767<=result767;
		result_out768<=result768;
		result_out769<=result769;
		result_out770<=result770;
		result_out771<=result771;
		result_out772<=result772;
		result_out773<=result773;
		result_out774<=result774;
		result_out775<=result775;
		result_out776<=result776;
		result_out777<=result777;
		result_out778<=result778;
		result_out779<=result779;
		result_out780<=result780;
		result_out781<=result781;
		result_out782<=result782;
		result_out783<=result783;
		result_out784<=result784;
		result_out785<=result785;
		result_out786<=result786;
		result_out787<=result787;
		result_out788<=result788;
		result_out789<=result789;
		result_out790<=result790;
		result_out791<=result791;
		result_out792<=result792;
		result_out793<=result793;
		result_out794<=result794;
		result_out795<=result795;
		result_out796<=result796;
		result_out797<=result797;
		result_out798<=result798;
		result_out799<=result799;
		result_out800<=result800;
		result_out801<=result801;
		result_out802<=result802;
		result_out803<=result803;
		result_out804<=result804;
		result_out805<=result805;
		result_out806<=result806;
		result_out807<=result807;
		result_out808<=result808;
		result_out809<=result809;
		result_out810<=result810;
		result_out811<=result811;
		result_out812<=result812;
		result_out813<=result813;
		result_out814<=result814;
		result_out815<=result815;
		result_out816<=result816;
		result_out817<=result817;
		result_out818<=result818;
		result_out819<=result819;
		result_out820<=result820;
		result_out821<=result821;
		result_out822<=result822;
		result_out823<=result823;
		result_out824<=result824;
		result_out825<=result825;
		result_out826<=result826;
		result_out827<=result827;
		result_out828<=result828;
		result_out829<=result829;
		result_out830<=result830;
		result_out831<=result831;
		result_out832<=result832;
		result_out833<=result833;
		result_out834<=result834;
		result_out835<=result835;
		result_out836<=result836;
		result_out837<=result837;
		result_out838<=result838;
		result_out839<=result839;
		result_out840<=result840;
		result_out841<=result841;
		result_out842<=result842;
		result_out843<=result843;
		result_out844<=result844;
		result_out845<=result845;
		result_out846<=result846;
		result_out847<=result847;
		result_out848<=result848;
		result_out849<=result849;
		result_out850<=result850;
		result_out851<=result851;
		result_out852<=result852;
		result_out853<=result853;
		result_out854<=result854;
		result_out855<=result855;
		result_out856<=result856;
		result_out857<=result857;
		result_out858<=result858;
		result_out859<=result859;
		result_out860<=result860;
		result_out861<=result861;
		result_out862<=result862;
		result_out863<=result863;
		result_out864<=result864;
		result_out865<=result865;
		result_out866<=result866;
		result_out867<=result867;
		result_out868<=result868;
		result_out869<=result869;
		result_out870<=result870;
		result_out871<=result871;
		result_out872<=result872;
		result_out873<=result873;
		result_out874<=result874;
		result_out875<=result875;
		result_out876<=result876;
		result_out877<=result877;
		result_out878<=result878;
		result_out879<=result879;
		result_out880<=result880;
		result_out881<=result881;
		result_out882<=result882;
		result_out883<=result883;
		result_out884<=result884;
		result_out885<=result885;
		result_out886<=result886;
		result_out887<=result887;
		result_out888<=result888;
		result_out889<=result889;
		result_out890<=result890;
		result_out891<=result891;
		result_out892<=result892;
		result_out893<=result893;
		result_out894<=result894;
		result_out895<=result895;
		result_out896<=result896;
		result_out897<=result897;
		result_out898<=result898;
		result_out899<=result899;
		result_out900<=result900;
		result_out901<=result901;
		result_out902<=result902;
		result_out903<=result903;
		result_out904<=result904;
		result_out905<=result905;
		result_out906<=result906;
		result_out907<=result907;
		result_out908<=result908;
		result_out909<=result909;
		result_out910<=result910;
		result_out911<=result911;
		result_out912<=result912;
		result_out913<=result913;
		result_out914<=result914;
		result_out915<=result915;
		result_out916<=result916;
		result_out917<=result917;
		result_out918<=result918;
		result_out919<=result919;
		result_out920<=result920;
		result_out921<=result921;
		result_out922<=result922;
		result_out923<=result923;
		result_out924<=result924;
		result_out925<=result925;
		result_out926<=result926;
		result_out927<=result927;
		result_out928<=result928;
		result_out929<=result929;
		result_out930<=result930;
		result_out931<=result931;
		result_out932<=result932;
		result_out933<=result933;
		result_out934<=result934;
		result_out935<=result935;
		result_out936<=result936;
		result_out937<=result937;
		result_out938<=result938;
		result_out939<=result939;
		result_out940<=result940;
		result_out941<=result941;
		result_out942<=result942;
		result_out943<=result943;
		result_out944<=result944;
		result_out945<=result945;
		result_out946<=result946;
		result_out947<=result947;
		result_out948<=result948;
		result_out949<=result949;
		result_out950<=result950;
		result_out951<=result951;
		result_out952<=result952;
		result_out953<=result953;
		result_out954<=result954;
		result_out955<=result955;
		result_out956<=result956;
		result_out957<=result957;
		result_out958<=result958;
		result_out959<=result959;
		result_out960<=result960;
		result_out961<=result961;
		result_out962<=result962;
		result_out963<=result963;
		result_out964<=result964;
		result_out965<=result965;
		result_out966<=result966;
		result_out967<=result967;
		result_out968<=result968;
		result_out969<=result969;
		result_out970<=result970;
		result_out971<=result971;
		result_out972<=result972;
		result_out973<=result973;
		result_out974<=result974;
		result_out975<=result975;
		result_out976<=result976;
		result_out977<=result977;
		result_out978<=result978;
		result_out979<=result979;
		result_out980<=result980;
		result_out981<=result981;
		result_out982<=result982;
		result_out983<=result983;
		result_out984<=result984;
		result_out985<=result985;
		result_out986<=result986;
		result_out987<=result987;
		result_out988<=result988;
		result_out989<=result989;
		result_out990<=result990;
		result_out991<=result991;
		result_out992<=result992;
		result_out993<=result993;
		result_out994<=result994;
		result_out995<=result995;
		result_out996<=result996;
		result_out997<=result997;
		result_out998<=result998;
		result_out999<=result999;
		result_out1000<=result1000;
		result_out1001<=result1001;
		result_out1002<=result1002;
		result_out1003<=result1003;
		result_out1004<=result1004;
		result_out1005<=result1005;
		result_out1006<=result1006;
		result_out1007<=result1007;
		result_out1008<=result1008;
		result_out1009<=result1009;
		result_out1010<=result1010;
		result_out1011<=result1011;
		result_out1012<=result1012;
		result_out1013<=result1013;
		result_out1014<=result1014;
		result_out1015<=result1015;
		result_out1016<=result1016;
		result_out1017<=result1017;
		result_out1018<=result1018;
		result_out1019<=result1019;
		result_out1020<=result1020;
		result_out1021<=result1021;
		result_out1022<=result1022;
		result_out1023<=result1023;
		result_out1024<=result1024;
		result_out1025<=result1025;
		result_out1026<=result1026;
		result_out1027<=result1027;
		result_out1028<=result1028;
		result_out1029<=result1029;
		result_out1030<=result1030;
		result_out1031<=result1031;
		result_out1032<=result1032;
		result_out1033<=result1033;
		result_out1034<=result1034;
		result_out1035<=result1035;
		result_out1036<=result1036;
		result_out1037<=result1037;
		result_out1038<=result1038;
		result_out1039<=result1039;
		result_out1040<=result1040;
		result_out1041<=result1041;
		result_out1042<=result1042;
		result_out1043<=result1043;
		result_out1044<=result1044;
		result_out1045<=result1045;
		result_out1046<=result1046;
		result_out1047<=result1047;
		result_out1048<=result1048;
		result_out1049<=result1049;
		result_out1050<=result1050;
		result_out1051<=result1051;
		result_out1052<=result1052;
		result_out1053<=result1053;
		result_out1054<=result1054;
		result_out1055<=result1055;
		result_out1056<=result1056;
		result_out1057<=result1057;
		result_out1058<=result1058;
		result_out1059<=result1059;
		result_out1060<=result1060;
		result_out1061<=result1061;
		result_out1062<=result1062;
		result_out1063<=result1063;
		result_out1064<=result1064;
		result_out1065<=result1065;
		result_out1066<=result1066;
		result_out1067<=result1067;
		result_out1068<=result1068;
		result_out1069<=result1069;
		result_out1070<=result1070;
		result_out1071<=result1071;
		result_out1072<=result1072;
		result_out1073<=result1073;
		result_out1074<=result1074;
		result_out1075<=result1075;
		result_out1076<=result1076;
		result_out1077<=result1077;
		result_out1078<=result1078;
		result_out1079<=result1079;
		result_out1080<=result1080;
		result_out1081<=result1081;
		result_out1082<=result1082;
		result_out1083<=result1083;
		result_out1084<=result1084;
		result_out1085<=result1085;
		result_out1086<=result1086;
		result_out1087<=result1087;
		result_out1088<=result1088;
		result_out1089<=result1089;
		result_out1090<=result1090;
		result_out1091<=result1091;
		result_out1092<=result1092;
		result_out1093<=result1093;
		result_out1094<=result1094;
		result_out1095<=result1095;
		result_out1096<=result1096;
		result_out1097<=result1097;
		result_out1098<=result1098;
		result_out1099<=result1099;
		result_out1100<=result1100;
		result_out1101<=result1101;
		result_out1102<=result1102;
		result_out1103<=result1103;
		result_out1104<=result1104;
		result_out1105<=result1105;
		result_out1106<=result1106;
		result_out1107<=result1107;
		result_out1108<=result1108;
		result_out1109<=result1109;
		result_out1110<=result1110;
		result_out1111<=result1111;
		result_out1112<=result1112;
		result_out1113<=result1113;
		result_out1114<=result1114;
		result_out1115<=result1115;
		result_out1116<=result1116;
		result_out1117<=result1117;
		result_out1118<=result1118;
		result_out1119<=result1119;
		result_out1120<=result1120;
		result_out1121<=result1121;
		result_out1122<=result1122;
		result_out1123<=result1123;
		result_out1124<=result1124;
		result_out1125<=result1125;
		result_out1126<=result1126;
		result_out1127<=result1127;
		result_out1128<=result1128;
		result_out1129<=result1129;
		result_out1130<=result1130;
		result_out1131<=result1131;
		result_out1132<=result1132;
		result_out1133<=result1133;
		result_out1134<=result1134;
		result_out1135<=result1135;
		result_out1136<=result1136;
		result_out1137<=result1137;
		result_out1138<=result1138;
		result_out1139<=result1139;
		result_out1140<=result1140;
		result_out1141<=result1141;
		result_out1142<=result1142;
		result_out1143<=result1143;
		result_out1144<=result1144;
		result_out1145<=result1145;
		result_out1146<=result1146;
		result_out1147<=result1147;
		result_out1148<=result1148;
		result_out1149<=result1149;
		result_out1150<=result1150;
		result_out1151<=result1151;
		result_out1152<=result1152;
		result_out1153<=result1153;
		result_out1154<=result1154;
		result_out1155<=result1155;
		result_out1156<=result1156;
		result_out1157<=result1157;
		result_out1158<=result1158;
		result_out1159<=result1159;
		result_out1160<=result1160;
		result_out1161<=result1161;
		result_out1162<=result1162;
		result_out1163<=result1163;
		result_out1164<=result1164;
		result_out1165<=result1165;
		result_out1166<=result1166;
		result_out1167<=result1167;
		result_out1168<=result1168;
		result_out1169<=result1169;
		result_out1170<=result1170;
		result_out1171<=result1171;
		result_out1172<=result1172;
		result_out1173<=result1173;
		result_out1174<=result1174;
		result_out1175<=result1175;
		result_out1176<=result1176;
		result_out1177<=result1177;
		result_out1178<=result1178;
		result_out1179<=result1179;
		result_out1180<=result1180;
		result_out1181<=result1181;
		result_out1182<=result1182;
		result_out1183<=result1183;
		result_out1184<=result1184;
		result_out1185<=result1185;
		result_out1186<=result1186;
		result_out1187<=result1187;
		result_out1188<=result1188;
		result_out1189<=result1189;
		result_out1190<=result1190;
		result_out1191<=result1191;
		result_out1192<=result1192;
		result_out1193<=result1193;
		result_out1194<=result1194;
		result_out1195<=result1195;
		result_out1196<=result1196;
		result_out1197<=result1197;
		result_out1198<=result1198;
		result_out1199<=result1199;
		result_out1200<=result1200;
		result_out1201<=result1201;
		result_out1202<=result1202;
		result_out1203<=result1203;
		result_out1204<=result1204;
		result_out1205<=result1205;
		result_out1206<=result1206;
		result_out1207<=result1207;
		result_out1208<=result1208;
		result_out1209<=result1209;
		result_out1210<=result1210;
		result_out1211<=result1211;
		result_out1212<=result1212;
		result_out1213<=result1213;
		result_out1214<=result1214;
		result_out1215<=result1215;
		result_out1216<=result1216;
		result_out1217<=result1217;
		result_out1218<=result1218;
		result_out1219<=result1219;
		result_out1220<=result1220;
		result_out1221<=result1221;
		result_out1222<=result1222;
		result_out1223<=result1223;
		result_out1224<=result1224;
		result_out1225<=result1225;
		result_out1226<=result1226;
		result_out1227<=result1227;
		result_out1228<=result1228;
		result_out1229<=result1229;
		result_out1230<=result1230;
		result_out1231<=result1231;
		result_out1232<=result1232;
		result_out1233<=result1233;
		result_out1234<=result1234;
		result_out1235<=result1235;
		result_out1236<=result1236;
		result_out1237<=result1237;
		result_out1238<=result1238;
		result_out1239<=result1239;
		result_out1240<=result1240;
		result_out1241<=result1241;
		result_out1242<=result1242;
		result_out1243<=result1243;
		result_out1244<=result1244;
		result_out1245<=result1245;
		result_out1246<=result1246;
		result_out1247<=result1247;
		result_out1248<=result1248;
		result_out1249<=result1249;
		result_out1250<=result1250;
		result_out1251<=result1251;
		result_out1252<=result1252;
		result_out1253<=result1253;
		result_out1254<=result1254;
		result_out1255<=result1255;
		result_out1256<=result1256;
		result_out1257<=result1257;
		result_out1258<=result1258;
		result_out1259<=result1259;
		result_out1260<=result1260;
		result_out1261<=result1261;
		result_out1262<=result1262;
		result_out1263<=result1263;
		result_out1264<=result1264;
		result_out1265<=result1265;
		result_out1266<=result1266;
		result_out1267<=result1267;
		result_out1268<=result1268;
		result_out1269<=result1269;
		result_out1270<=result1270;
		result_out1271<=result1271;
		result_out1272<=result1272;
		result_out1273<=result1273;
		result_out1274<=result1274;
		result_out1275<=result1275;
		result_out1276<=result1276;
		result_out1277<=result1277;
		result_out1278<=result1278;
		result_out1279<=result1279;
		result_out1280<=result1280;
		result_out1281<=result1281;
		result_out1282<=result1282;
		result_out1283<=result1283;
		result_out1284<=result1284;
		result_out1285<=result1285;
		result_out1286<=result1286;
		result_out1287<=result1287;
		result_out1288<=result1288;
		result_out1289<=result1289;
		result_out1290<=result1290;
		result_out1291<=result1291;
		result_out1292<=result1292;
		result_out1293<=result1293;
		result_out1294<=result1294;
		result_out1295<=result1295;
		result_out1296<=result1296;
		result_out1297<=result1297;
		result_out1298<=result1298;
		result_out1299<=result1299;
		result_out1300<=result1300;
		result_out1301<=result1301;
		result_out1302<=result1302;
		result_out1303<=result1303;
		result_out1304<=result1304;
		result_out1305<=result1305;
		result_out1306<=result1306;
		result_out1307<=result1307;
		result_out1308<=result1308;
		result_out1309<=result1309;
		result_out1310<=result1310;
		result_out1311<=result1311;
		result_out1312<=result1312;
		result_out1313<=result1313;
		result_out1314<=result1314;
		result_out1315<=result1315;
		result_out1316<=result1316;
		result_out1317<=result1317;
		result_out1318<=result1318;
		result_out1319<=result1319;
		result_out1320<=result1320;
		result_out1321<=result1321;
		result_out1322<=result1322;
		result_out1323<=result1323;
		result_out1324<=result1324;
		result_out1325<=result1325;
		result_out1326<=result1326;
		result_out1327<=result1327;
		result_out1328<=result1328;
		result_out1329<=result1329;
		result_out1330<=result1330;
		result_out1331<=result1331;
		result_out1332<=result1332;
		result_out1333<=result1333;
		result_out1334<=result1334;
		result_out1335<=result1335;
		result_out1336<=result1336;
		result_out1337<=result1337;
		result_out1338<=result1338;
		result_out1339<=result1339;
		result_out1340<=result1340;
		result_out1341<=result1341;
		result_out1342<=result1342;
		result_out1343<=result1343;
		result_out1344<=result1344;
		result_out1345<=result1345;
		result_out1346<=result1346;
		result_out1347<=result1347;
		result_out1348<=result1348;
		result_out1349<=result1349;
		result_out1350<=result1350;
		result_out1351<=result1351;
		result_out1352<=result1352;
		result_out1353<=result1353;
		result_out1354<=result1354;
		result_out1355<=result1355;
		result_out1356<=result1356;
		result_out1357<=result1357;
		result_out1358<=result1358;
		result_out1359<=result1359;
		result_out1360<=result1360;
		result_out1361<=result1361;
		result_out1362<=result1362;
		result_out1363<=result1363;
		result_out1364<=result1364;
		result_out1365<=result1365;
		result_out1366<=result1366;
		result_out1367<=result1367;
		result_out1368<=result1368;
		result_out1369<=result1369;
		result_out1370<=result1370;
		result_out1371<=result1371;
		result_out1372<=result1372;
		result_out1373<=result1373;
		result_out1374<=result1374;
		result_out1375<=result1375;
		result_out1376<=result1376;
		result_out1377<=result1377;
		result_out1378<=result1378;
		result_out1379<=result1379;
		result_out1380<=result1380;
		result_out1381<=result1381;
		result_out1382<=result1382;
		result_out1383<=result1383;
		result_out1384<=result1384;
		result_out1385<=result1385;
		result_out1386<=result1386;
		result_out1387<=result1387;
		result_out1388<=result1388;
		result_out1389<=result1389;
		result_out1390<=result1390;
		result_out1391<=result1391;
		result_out1392<=result1392;
		result_out1393<=result1393;
		result_out1394<=result1394;
		result_out1395<=result1395;
		result_out1396<=result1396;
		result_out1397<=result1397;
		result_out1398<=result1398;
		result_out1399<=result1399;
		result_out1400<=result1400;
		result_out1401<=result1401;
		result_out1402<=result1402;
		result_out1403<=result1403;
		result_out1404<=result1404;
		result_out1405<=result1405;
		result_out1406<=result1406;
		result_out1407<=result1407;
		result_out1408<=result1408;
		result_out1409<=result1409;
		result_out1410<=result1410;
		result_out1411<=result1411;
		result_out1412<=result1412;
		result_out1413<=result1413;
		result_out1414<=result1414;
		result_out1415<=result1415;
		result_out1416<=result1416;
		result_out1417<=result1417;
		result_out1418<=result1418;
		result_out1419<=result1419;
		result_out1420<=result1420;
		result_out1421<=result1421;
		result_out1422<=result1422;
		result_out1423<=result1423;
		result_out1424<=result1424;
		result_out1425<=result1425;
		result_out1426<=result1426;
		result_out1427<=result1427;
		result_out1428<=result1428;
		result_out1429<=result1429;
		result_out1430<=result1430;
		result_out1431<=result1431;
		result_out1432<=result1432;
		result_out1433<=result1433;
		result_out1434<=result1434;
		result_out1435<=result1435;
		result_out1436<=result1436;
		result_out1437<=result1437;
		result_out1438<=result1438;
		result_out1439<=result1439;
		result_out1440<=result1440;
		result_out1441<=result1441;
		result_out1442<=result1442;
		result_out1443<=result1443;
		result_out1444<=result1444;
		result_out1445<=result1445;
		result_out1446<=result1446;
		result_out1447<=result1447;
		result_out1448<=result1448;
		result_out1449<=result1449;
		result_out1450<=result1450;
		result_out1451<=result1451;
		result_out1452<=result1452;
		result_out1453<=result1453;
		result_out1454<=result1454;
		result_out1455<=result1455;
		result_out1456<=result1456;
		result_out1457<=result1457;
		result_out1458<=result1458;
		result_out1459<=result1459;
		result_out1460<=result1460;
		result_out1461<=result1461;
		result_out1462<=result1462;
		result_out1463<=result1463;
		result_out1464<=result1464;
		result_out1465<=result1465;
		result_out1466<=result1466;
		result_out1467<=result1467;
		result_out1468<=result1468;
		result_out1469<=result1469;
		result_out1470<=result1470;
		result_out1471<=result1471;
		result_out1472<=result1472;
		result_out1473<=result1473;
		result_out1474<=result1474;
		result_out1475<=result1475;
		result_out1476<=result1476;
		result_out1477<=result1477;
		result_out1478<=result1478;
		result_out1479<=result1479;
		result_out1480<=result1480;
		result_out1481<=result1481;
		result_out1482<=result1482;
		result_out1483<=result1483;
		result_out1484<=result1484;
		result_out1485<=result1485;
		result_out1486<=result1486;
		result_out1487<=result1487;
		result_out1488<=result1488;
		result_out1489<=result1489;
		result_out1490<=result1490;
		result_out1491<=result1491;
		result_out1492<=result1492;
		result_out1493<=result1493;
		result_out1494<=result1494;
		result_out1495<=result1495;
		result_out1496<=result1496;
		result_out1497<=result1497;
		result_out1498<=result1498;
		result_out1499<=result1499;
		result_out1500<=result1500;
		result_out1501<=result1501;
		result_out1502<=result1502;
		result_out1503<=result1503;
		result_out1504<=result1504;
		result_out1505<=result1505;
		result_out1506<=result1506;
		result_out1507<=result1507;
		result_out1508<=result1508;
		result_out1509<=result1509;
		result_out1510<=result1510;
		result_out1511<=result1511;
		result_out1512<=result1512;
		result_out1513<=result1513;
		result_out1514<=result1514;
		result_out1515<=result1515;
		result_out1516<=result1516;
		result_out1517<=result1517;
		result_out1518<=result1518;
		result_out1519<=result1519;
		result_out1520<=result1520;
		result_out1521<=result1521;
		result_out1522<=result1522;
		result_out1523<=result1523;
		result_out1524<=result1524;
		result_out1525<=result1525;
		result_out1526<=result1526;
		result_out1527<=result1527;
		result_out1528<=result1528;
		result_out1529<=result1529;
		result_out1530<=result1530;
		result_out1531<=result1531;
		result_out1532<=result1532;
		result_out1533<=result1533;
		result_out1534<=result1534;
		result_out1535<=result1535;
		result_out1536<=result1536;
		result_out1537<=result1537;
		result_out1538<=result1538;
		result_out1539<=result1539;
		result_out1540<=result1540;
		result_out1541<=result1541;
		result_out1542<=result1542;
		result_out1543<=result1543;
		result_out1544<=result1544;
		result_out1545<=result1545;
		result_out1546<=result1546;
		result_out1547<=result1547;
		result_out1548<=result1548;
		result_out1549<=result1549;
		result_out1550<=result1550;
		result_out1551<=result1551;
		result_out1552<=result1552;
		result_out1553<=result1553;
		result_out1554<=result1554;
		result_out1555<=result1555;
		result_out1556<=result1556;
		result_out1557<=result1557;
		result_out1558<=result1558;
		result_out1559<=result1559;
		result_out1560<=result1560;
		result_out1561<=result1561;
		result_out1562<=result1562;
		result_out1563<=result1563;
		result_out1564<=result1564;
		result_out1565<=result1565;
		result_out1566<=result1566;
		result_out1567<=result1567;
		result_out1568<=result1568;
		result_out1569<=result1569;
		result_out1570<=result1570;
		result_out1571<=result1571;
		result_out1572<=result1572;
		result_out1573<=result1573;
		result_out1574<=result1574;
		result_out1575<=result1575;
		result_out1576<=result1576;
		result_out1577<=result1577;
		result_out1578<=result1578;
		result_out1579<=result1579;
		result_out1580<=result1580;
		result_out1581<=result1581;
		result_out1582<=result1582;
		result_out1583<=result1583;
		result_out1584<=result1584;
		result_out1585<=result1585;
		result_out1586<=result1586;
		result_out1587<=result1587;
		result_out1588<=result1588;
		result_out1589<=result1589;
		result_out1590<=result1590;
		result_out1591<=result1591;
		result_out1592<=result1592;
		result_out1593<=result1593;
		result_out1594<=result1594;
		result_out1595<=result1595;
		result_out1596<=result1596;
		result_out1597<=result1597;
		result_out1598<=result1598;
		result_out1599<=result1599;
		result_out1600<=result1600;
		result_out1601<=result1601;
		result_out1602<=result1602;
		result_out1603<=result1603;
		result_out1604<=result1604;
		result_out1605<=result1605;
		result_out1606<=result1606;
		result_out1607<=result1607;
		result_out1608<=result1608;
		result_out1609<=result1609;
		result_out1610<=result1610;
		result_out1611<=result1611;
		result_out1612<=result1612;
		result_out1613<=result1613;
		result_out1614<=result1614;
		result_out1615<=result1615;
		result_out1616<=result1616;
		result_out1617<=result1617;
		result_out1618<=result1618;
		result_out1619<=result1619;
		result_out1620<=result1620;
		result_out1621<=result1621;
		result_out1622<=result1622;
		result_out1623<=result1623;
		result_out1624<=result1624;
		result_out1625<=result1625;
		result_out1626<=result1626;
		result_out1627<=result1627;
		result_out1628<=result1628;
		result_out1629<=result1629;
		result_out1630<=result1630;
		result_out1631<=result1631;
		result_out1632<=result1632;
		result_out1633<=result1633;
		result_out1634<=result1634;
		result_out1635<=result1635;
		result_out1636<=result1636;
		result_out1637<=result1637;
		result_out1638<=result1638;
		result_out1639<=result1639;
		result_out1640<=result1640;
		result_out1641<=result1641;
		result_out1642<=result1642;
		result_out1643<=result1643;
		result_out1644<=result1644;
		result_out1645<=result1645;
		result_out1646<=result1646;
		result_out1647<=result1647;
		result_out1648<=result1648;
		result_out1649<=result1649;
		result_out1650<=result1650;
		result_out1651<=result1651;
		result_out1652<=result1652;
		result_out1653<=result1653;
		result_out1654<=result1654;
		result_out1655<=result1655;
		result_out1656<=result1656;
		result_out1657<=result1657;
		result_out1658<=result1658;
		result_out1659<=result1659;
		result_out1660<=result1660;
		result_out1661<=result1661;
		result_out1662<=result1662;
		result_out1663<=result1663;
		result_out1664<=result1664;
		result_out1665<=result1665;
		result_out1666<=result1666;
		result_out1667<=result1667;
		result_out1668<=result1668;
		result_out1669<=result1669;
		result_out1670<=result1670;
		result_out1671<=result1671;
		result_out1672<=result1672;
		result_out1673<=result1673;
		result_out1674<=result1674;
		result_out1675<=result1675;
		result_out1676<=result1676;
		result_out1677<=result1677;
		result_out1678<=result1678;
		result_out1679<=result1679;
		result_out1680<=result1680;
		result_out1681<=result1681;
		result_out1682<=result1682;
		result_out1683<=result1683;
		result_out1684<=result1684;
		result_out1685<=result1685;
		result_out1686<=result1686;
		result_out1687<=result1687;
		result_out1688<=result1688;
		result_out1689<=result1689;
		result_out1690<=result1690;
		result_out1691<=result1691;
		result_out1692<=result1692;
		result_out1693<=result1693;
		result_out1694<=result1694;
		result_out1695<=result1695;
		result_out1696<=result1696;
		result_out1697<=result1697;
		result_out1698<=result1698;
		result_out1699<=result1699;
		result_out1700<=result1700;
		result_out1701<=result1701;
		result_out1702<=result1702;
		result_out1703<=result1703;
		result_out1704<=result1704;
		result_out1705<=result1705;
		result_out1706<=result1706;
		result_out1707<=result1707;
		result_out1708<=result1708;
		result_out1709<=result1709;
		result_out1710<=result1710;
		result_out1711<=result1711;
		result_out1712<=result1712;
		result_out1713<=result1713;
		result_out1714<=result1714;
		result_out1715<=result1715;
		result_out1716<=result1716;
		result_out1717<=result1717;
		result_out1718<=result1718;
		result_out1719<=result1719;
		result_out1720<=result1720;
		result_out1721<=result1721;
		result_out1722<=result1722;
		result_out1723<=result1723;
		result_out1724<=result1724;
		result_out1725<=result1725;
		result_out1726<=result1726;
		result_out1727<=result1727;
		result_out1728<=result1728;
		result_out1729<=result1729;
		result_out1730<=result1730;
		result_out1731<=result1731;
		result_out1732<=result1732;
		result_out1733<=result1733;
		result_out1734<=result1734;
		result_out1735<=result1735;
		result_out1736<=result1736;
		result_out1737<=result1737;
		result_out1738<=result1738;
		result_out1739<=result1739;
		result_out1740<=result1740;
		result_out1741<=result1741;
		result_out1742<=result1742;
		result_out1743<=result1743;
		result_out1744<=result1744;
		result_out1745<=result1745;
		result_out1746<=result1746;
		result_out1747<=result1747;
		result_out1748<=result1748;
		result_out1749<=result1749;
		result_out1750<=result1750;
		result_out1751<=result1751;
		result_out1752<=result1752;
		result_out1753<=result1753;
		result_out1754<=result1754;
		result_out1755<=result1755;
		result_out1756<=result1756;
		result_out1757<=result1757;
		result_out1758<=result1758;
		result_out1759<=result1759;
		result_out1760<=result1760;
		result_out1761<=result1761;
		result_out1762<=result1762;
		result_out1763<=result1763;
		result_out1764<=result1764;
		result_out1765<=result1765;
		result_out1766<=result1766;
		result_out1767<=result1767;
		result_out1768<=result1768;
		result_out1769<=result1769;
		result_out1770<=result1770;
		result_out1771<=result1771;
		result_out1772<=result1772;
		result_out1773<=result1773;
		result_out1774<=result1774;
		result_out1775<=result1775;
		result_out1776<=result1776;
		result_out1777<=result1777;
		result_out1778<=result1778;
		result_out1779<=result1779;
		result_out1780<=result1780;
		result_out1781<=result1781;
		result_out1782<=result1782;
		result_out1783<=result1783;
		result_out1784<=result1784;
		result_out1785<=result1785;
		result_out1786<=result1786;
		result_out1787<=result1787;
		result_out1788<=result1788;
		result_out1789<=result1789;
		result_out1790<=result1790;
		result_out1791<=result1791;
		result_out1792<=result1792;
		result_out1793<=result1793;
		result_out1794<=result1794;
		result_out1795<=result1795;
		result_out1796<=result1796;
		result_out1797<=result1797;
		result_out1798<=result1798;
		result_out1799<=result1799;
		result_out1800<=result1800;
		result_out1801<=result1801;
		result_out1802<=result1802;
		result_out1803<=result1803;
		result_out1804<=result1804;
		result_out1805<=result1805;
		result_out1806<=result1806;
		result_out1807<=result1807;
		result_out1808<=result1808;
		result_out1809<=result1809;
		result_out1810<=result1810;
		result_out1811<=result1811;
		result_out1812<=result1812;
		result_out1813<=result1813;
		result_out1814<=result1814;
		result_out1815<=result1815;
		result_out1816<=result1816;
		result_out1817<=result1817;
		result_out1818<=result1818;
		result_out1819<=result1819;
		result_out1820<=result1820;
		result_out1821<=result1821;
		result_out1822<=result1822;
		result_out1823<=result1823;
		result_out1824<=result1824;
		result_out1825<=result1825;
		result_out1826<=result1826;
		result_out1827<=result1827;
		result_out1828<=result1828;
		result_out1829<=result1829;
		result_out1830<=result1830;
		result_out1831<=result1831;
		result_out1832<=result1832;
		result_out1833<=result1833;
		result_out1834<=result1834;
		result_out1835<=result1835;
		result_out1836<=result1836;
		result_out1837<=result1837;
		result_out1838<=result1838;
		result_out1839<=result1839;
		result_out1840<=result1840;
		result_out1841<=result1841;
		result_out1842<=result1842;
		result_out1843<=result1843;
		result_out1844<=result1844;
		result_out1845<=result1845;
		result_out1846<=result1846;
		result_out1847<=result1847;
		result_out1848<=result1848;
		result_out1849<=result1849;
		result_out1850<=result1850;
		result_out1851<=result1851;
		result_out1852<=result1852;
		result_out1853<=result1853;
		result_out1854<=result1854;
		result_out1855<=result1855;
		result_out1856<=result1856;
		result_out1857<=result1857;
		result_out1858<=result1858;
		result_out1859<=result1859;
		result_out1860<=result1860;
		result_out1861<=result1861;
		result_out1862<=result1862;
		result_out1863<=result1863;
		result_out1864<=result1864;
		result_out1865<=result1865;
		result_out1866<=result1866;
		result_out1867<=result1867;
		result_out1868<=result1868;
		result_out1869<=result1869;
		result_out1870<=result1870;
		result_out1871<=result1871;
		result_out1872<=result1872;
		result_out1873<=result1873;
		result_out1874<=result1874;
		result_out1875<=result1875;
		result_out1876<=result1876;
		result_out1877<=result1877;
		result_out1878<=result1878;
		result_out1879<=result1879;
		result_out1880<=result1880;
		result_out1881<=result1881;
		result_out1882<=result1882;
		result_out1883<=result1883;
		result_out1884<=result1884;
		result_out1885<=result1885;
		result_out1886<=result1886;
		result_out1887<=result1887;
		result_out1888<=result1888;
		result_out1889<=result1889;
		result_out1890<=result1890;
		result_out1891<=result1891;
		result_out1892<=result1892;
		result_out1893<=result1893;
		result_out1894<=result1894;
		result_out1895<=result1895;
		result_out1896<=result1896;
		result_out1897<=result1897;
		result_out1898<=result1898;
		result_out1899<=result1899;
		result_out1900<=result1900;
		result_out1901<=result1901;
		result_out1902<=result1902;
		result_out1903<=result1903;
		result_out1904<=result1904;
		result_out1905<=result1905;
		result_out1906<=result1906;
		result_out1907<=result1907;
		result_out1908<=result1908;
		result_out1909<=result1909;
		result_out1910<=result1910;
		result_out1911<=result1911;
		result_out1912<=result1912;
		result_out1913<=result1913;
		result_out1914<=result1914;
		result_out1915<=result1915;
		result_out1916<=result1916;
		result_out1917<=result1917;
		result_out1918<=result1918;
		result_out1919<=result1919;
		result_out1920<=result1920;
		result_out1921<=result1921;
		result_out1922<=result1922;
		result_out1923<=result1923;
		result_out1924<=result1924;
		result_out1925<=result1925;
		result_out1926<=result1926;
		result_out1927<=result1927;
		result_out1928<=result1928;
		result_out1929<=result1929;
		result_out1930<=result1930;
		result_out1931<=result1931;
		result_out1932<=result1932;
		result_out1933<=result1933;
		result_out1934<=result1934;
		result_out1935<=result1935;
		result_out1936<=result1936;
		result_out1937<=result1937;
		result_out1938<=result1938;
		result_out1939<=result1939;
		result_out1940<=result1940;
		result_out1941<=result1941;
		result_out1942<=result1942;
		result_out1943<=result1943;
		result_out1944<=result1944;
		result_out1945<=result1945;
		result_out1946<=result1946;
		result_out1947<=result1947;
		result_out1948<=result1948;
		result_out1949<=result1949;
		result_out1950<=result1950;
		result_out1951<=result1951;
		result_out1952<=result1952;
		result_out1953<=result1953;
		result_out1954<=result1954;
		result_out1955<=result1955;
		result_out1956<=result1956;
		result_out1957<=result1957;
		result_out1958<=result1958;
		result_out1959<=result1959;
		result_out1960<=result1960;
		result_out1961<=result1961;
		result_out1962<=result1962;
		result_out1963<=result1963;
		result_out1964<=result1964;
		result_out1965<=result1965;
		result_out1966<=result1966;
		result_out1967<=result1967;
		result_out1968<=result1968;
		result_out1969<=result1969;
		result_out1970<=result1970;
		result_out1971<=result1971;
		result_out1972<=result1972;
		result_out1973<=result1973;
		result_out1974<=result1974;
		result_out1975<=result1975;
		result_out1976<=result1976;
		result_out1977<=result1977;
		result_out1978<=result1978;
		result_out1979<=result1979;
		result_out1980<=result1980;
		result_out1981<=result1981;
		result_out1982<=result1982;
		result_out1983<=result1983;
		result_out1984<=result1984;
		result_out1985<=result1985;
		result_out1986<=result1986;
		result_out1987<=result1987;
		result_out1988<=result1988;
		result_out1989<=result1989;
		result_out1990<=result1990;
		result_out1991<=result1991;
		result_out1992<=result1992;
		result_out1993<=result1993;
		result_out1994<=result1994;
		result_out1995<=result1995;
		result_out1996<=result1996;
		result_out1997<=result1997;
		result_out1998<=result1998;
		result_out1999<=result1999;
		result_out2000<=result2000;
		result_out2001<=result2001;
		result_out2002<=result2002;
		result_out2003<=result2003;
		result_out2004<=result2004;
		result_out2005<=result2005;
		result_out2006<=result2006;
		result_out2007<=result2007;
		result_out2008<=result2008;
		result_out2009<=result2009;
		result_out2010<=result2010;
		result_out2011<=result2011;
		result_out2012<=result2012;
		result_out2013<=result2013;
		result_out2014<=result2014;
		result_out2015<=result2015;
		result_out2016<=result2016;
		result_out2017<=result2017;
		result_out2018<=result2018;
		result_out2019<=result2019;
		result_out2020<=result2020;
		result_out2021<=result2021;
		result_out2022<=result2022;
		result_out2023<=result2023;
		result_out2024<=result2024;
		result_out2025<=result2025;
		result_out2026<=result2026;
		result_out2027<=result2027;
		result_out2028<=result2028;
		result_out2029<=result2029;
		result_out2030<=result2030;
		result_out2031<=result2031;
		result_out2032<=result2032;
		result_out2033<=result2033;
		result_out2034<=result2034;
		result_out2035<=result2035;
		result_out2036<=result2036;
		result_out2037<=result2037;
		result_out2038<=result2038;
		result_out2039<=result2039;
		result_out2040<=result2040;
		result_out2041<=result2041;
		result_out2042<=result2042;
		result_out2043<=result2043;
		result_out2044<=result2044;
		result_out2045<=result2045;
		result_out2046<=result2046;
		result_out2047<=result2047;
		result_out2048<=result2048;
		result_out2049<=result2049;
		result_out2050<=result2050;
		result_out2051<=result2051;
		result_out2052<=result2052;
		result_out2053<=result2053;
		result_out2054<=result2054;
		result_out2055<=result2055;
		result_out2056<=result2056;
		result_out2057<=result2057;
		result_out2058<=result2058;
		result_out2059<=result2059;
		result_out2060<=result2060;
		result_out2061<=result2061;
		result_out2062<=result2062;
		result_out2063<=result2063;
		result_out2064<=result2064;
		result_out2065<=result2065;
		result_out2066<=result2066;
		result_out2067<=result2067;
		result_out2068<=result2068;
		result_out2069<=result2069;
		result_out2070<=result2070;
		result_out2071<=result2071;
		result_out2072<=result2072;
		result_out2073<=result2073;
		result_out2074<=result2074;
		result_out2075<=result2075;
		result_out2076<=result2076;
		result_out2077<=result2077;
		result_out2078<=result2078;
		result_out2079<=result2079;
		result_out2080<=result2080;
		result_out2081<=result2081;
		result_out2082<=result2082;
		result_out2083<=result2083;
		result_out2084<=result2084;
		result_out2085<=result2085;
		result_out2086<=result2086;
		result_out2087<=result2087;
		result_out2088<=result2088;
		result_out2089<=result2089;
		result_out2090<=result2090;
		result_out2091<=result2091;
		result_out2092<=result2092;
		result_out2093<=result2093;
		result_out2094<=result2094;
		result_out2095<=result2095;
		result_out2096<=result2096;
		result_out2097<=result2097;
		result_out2098<=result2098;
		result_out2099<=result2099;
		result_out2100<=result2100;
		result_out2101<=result2101;
		result_out2102<=result2102;
		result_out2103<=result2103;
		result_out2104<=result2104;
		result_out2105<=result2105;
		result_out2106<=result2106;
		result_out2107<=result2107;
		result_out2108<=result2108;
		result_out2109<=result2109;
		result_out2110<=result2110;
		result_out2111<=result2111;
		result_out2112<=result2112;
		result_out2113<=result2113;
		result_out2114<=result2114;
		result_out2115<=result2115;
		result_out2116<=result2116;
		result_out2117<=result2117;
		result_out2118<=result2118;
		result_out2119<=result2119;
		result_out2120<=result2120;
		result_out2121<=result2121;
		result_out2122<=result2122;
		result_out2123<=result2123;
		result_out2124<=result2124;
		result_out2125<=result2125;
		result_out2126<=result2126;
		result_out2127<=result2127;
		result_out2128<=result2128;
		result_out2129<=result2129;
		result_out2130<=result2130;
		result_out2131<=result2131;
		result_out2132<=result2132;
		result_out2133<=result2133;
		result_out2134<=result2134;
		result_out2135<=result2135;
		result_out2136<=result2136;
		result_out2137<=result2137;
		result_out2138<=result2138;
		result_out2139<=result2139;
		result_out2140<=result2140;
		result_out2141<=result2141;
		result_out2142<=result2142;
		result_out2143<=result2143;
		result_out2144<=result2144;
		result_out2145<=result2145;
		result_out2146<=result2146;
		result_out2147<=result2147;
		result_out2148<=result2148;
		result_out2149<=result2149;
		result_out2150<=result2150;
		result_out2151<=result2151;
		result_out2152<=result2152;
		result_out2153<=result2153;
		result_out2154<=result2154;
		result_out2155<=result2155;
		result_out2156<=result2156;
		result_out2157<=result2157;
		result_out2158<=result2158;
		result_out2159<=result2159;
		result_out2160<=result2160;
		result_out2161<=result2161;
		result_out2162<=result2162;
		result_out2163<=result2163;
		result_out2164<=result2164;
		result_out2165<=result2165;
		result_out2166<=result2166;
		result_out2167<=result2167;
		result_out2168<=result2168;
		result_out2169<=result2169;
		result_out2170<=result2170;
		result_out2171<=result2171;
		result_out2172<=result2172;
		result_out2173<=result2173;
		result_out2174<=result2174;
		result_out2175<=result2175;
		result_out2176<=result2176;
		result_out2177<=result2177;
		result_out2178<=result2178;
		result_out2179<=result2179;
		result_out2180<=result2180;
		result_out2181<=result2181;
		result_out2182<=result2182;
		result_out2183<=result2183;
		result_out2184<=result2184;
		result_out2185<=result2185;
		result_out2186<=result2186;
		result_out2187<=result2187;
		result_out2188<=result2188;
		result_out2189<=result2189;
		result_out2190<=result2190;
		result_out2191<=result2191;
		result_out2192<=result2192;
		result_out2193<=result2193;
		result_out2194<=result2194;
		result_out2195<=result2195;
		result_out2196<=result2196;
		result_out2197<=result2197;
		result_out2198<=result2198;
		result_out2199<=result2199;
		result_out2200<=result2200;
		result_out2201<=result2201;
		result_out2202<=result2202;
		result_out2203<=result2203;
		result_out2204<=result2204;
		result_out2205<=result2205;
		result_out2206<=result2206;
		result_out2207<=result2207;
		result_out2208<=result2208;
		result_out2209<=result2209;
		result_out2210<=result2210;
		result_out2211<=result2211;
		result_out2212<=result2212;
		result_out2213<=result2213;
		result_out2214<=result2214;
		result_out2215<=result2215;
		result_out2216<=result2216;
		result_out2217<=result2217;
		result_out2218<=result2218;
		result_out2219<=result2219;
		result_out2220<=result2220;
		result_out2221<=result2221;
		result_out2222<=result2222;
		result_out2223<=result2223;
		result_out2224<=result2224;
		result_out2225<=result2225;
		result_out2226<=result2226;
		result_out2227<=result2227;
		result_out2228<=result2228;
		result_out2229<=result2229;
		result_out2230<=result2230;
		result_out2231<=result2231;
		result_out2232<=result2232;
		result_out2233<=result2233;
		result_out2234<=result2234;
		result_out2235<=result2235;
		result_out2236<=result2236;
		result_out2237<=result2237;
		result_out2238<=result2238;
		result_out2239<=result2239;
		result_out2240<=result2240;
		result_out2241<=result2241;
		result_out2242<=result2242;
		result_out2243<=result2243;
		result_out2244<=result2244;
		result_out2245<=result2245;
		result_out2246<=result2246;
		result_out2247<=result2247;
		result_out2248<=result2248;
		result_out2249<=result2249;
		result_out2250<=result2250;
		result_out2251<=result2251;
		result_out2252<=result2252;
		result_out2253<=result2253;
		result_out2254<=result2254;
		result_out2255<=result2255;
		result_out2256<=result2256;
		result_out2257<=result2257;
		result_out2258<=result2258;
		result_out2259<=result2259;
		result_out2260<=result2260;
		result_out2261<=result2261;
		result_out2262<=result2262;
		result_out2263<=result2263;
		result_out2264<=result2264;
		result_out2265<=result2265;
		result_out2266<=result2266;
		result_out2267<=result2267;
		result_out2268<=result2268;
		result_out2269<=result2269;
		result_out2270<=result2270;
		result_out2271<=result2271;
		result_out2272<=result2272;
		result_out2273<=result2273;
		result_out2274<=result2274;
		result_out2275<=result2275;
		result_out2276<=result2276;
		result_out2277<=result2277;
		result_out2278<=result2278;
		result_out2279<=result2279;
		result_out2280<=result2280;
		result_out2281<=result2281;
		result_out2282<=result2282;
		result_out2283<=result2283;
		result_out2284<=result2284;
		result_out2285<=result2285;
		result_out2286<=result2286;
		result_out2287<=result2287;
		result_out2288<=result2288;
		result_out2289<=result2289;
		result_out2290<=result2290;
		result_out2291<=result2291;
		result_out2292<=result2292;
		result_out2293<=result2293;
		result_out2294<=result2294;
		result_out2295<=result2295;
		result_out2296<=result2296;
		result_out2297<=result2297;
		result_out2298<=result2298;
		result_out2299<=result2299;
		result_out2300<=result2300;
		result_out2301<=result2301;
		result_out2302<=result2302;
		result_out2303<=result2303;
		result_out2304<=result2304;
		result_out2305<=result2305;
		result_out2306<=result2306;
		result_out2307<=result2307;
		result_out2308<=result2308;
		result_out2309<=result2309;
		result_out2310<=result2310;
		result_out2311<=result2311;
		result_out2312<=result2312;
		result_out2313<=result2313;
		result_out2314<=result2314;
		result_out2315<=result2315;
		result_out2316<=result2316;
		result_out2317<=result2317;
		result_out2318<=result2318;
		result_out2319<=result2319;
		result_out2320<=result2320;
		result_out2321<=result2321;
		result_out2322<=result2322;
		result_out2323<=result2323;
		result_out2324<=result2324;
		result_out2325<=result2325;
		result_out2326<=result2326;
		result_out2327<=result2327;
		result_out2328<=result2328;
		result_out2329<=result2329;
		result_out2330<=result2330;
		result_out2331<=result2331;
		result_out2332<=result2332;
		result_out2333<=result2333;
		result_out2334<=result2334;
		result_out2335<=result2335;
		result_out2336<=result2336;
		result_out2337<=result2337;
		result_out2338<=result2338;
		result_out2339<=result2339;
		result_out2340<=result2340;
		result_out2341<=result2341;
		result_out2342<=result2342;
		result_out2343<=result2343;
		result_out2344<=result2344;
		result_out2345<=result2345;
		result_out2346<=result2346;
		result_out2347<=result2347;
		result_out2348<=result2348;
		result_out2349<=result2349;
		result_out2350<=result2350;
		result_out2351<=result2351;
		result_out2352<=result2352;
		result_out2353<=result2353;
		result_out2354<=result2354;
		result_out2355<=result2355;
		result_out2356<=result2356;
		result_out2357<=result2357;
		result_out2358<=result2358;
		result_out2359<=result2359;
		result_out2360<=result2360;
		result_out2361<=result2361;
		result_out2362<=result2362;
		result_out2363<=result2363;
		result_out2364<=result2364;
		result_out2365<=result2365;
		result_out2366<=result2366;
		result_out2367<=result2367;
		result_out2368<=result2368;
		result_out2369<=result2369;
		result_out2370<=result2370;
		result_out2371<=result2371;
		result_out2372<=result2372;
		result_out2373<=result2373;
		result_out2374<=result2374;
		result_out2375<=result2375;
		result_out2376<=result2376;
		result_out2377<=result2377;
		result_out2378<=result2378;
		result_out2379<=result2379;
		result_out2380<=result2380;
		result_out2381<=result2381;
		result_out2382<=result2382;
		result_out2383<=result2383;
		result_out2384<=result2384;
		result_out2385<=result2385;
		result_out2386<=result2386;
		result_out2387<=result2387;
		result_out2388<=result2388;
		result_out2389<=result2389;
		result_out2390<=result2390;
		result_out2391<=result2391;
		result_out2392<=result2392;
		result_out2393<=result2393;
		result_out2394<=result2394;
		result_out2395<=result2395;
		result_out2396<=result2396;
		result_out2397<=result2397;
		result_out2398<=result2398;
		result_out2399<=result2399;
		result_out2400<=result2400;
		result_out2401<=result2401;
		result_out2402<=result2402;
		result_out2403<=result2403;
		result_out2404<=result2404;
		result_out2405<=result2405;
		result_out2406<=result2406;
		result_out2407<=result2407;
		result_out2408<=result2408;
		result_out2409<=result2409;
		result_out2410<=result2410;
		result_out2411<=result2411;
		result_out2412<=result2412;
		result_out2413<=result2413;
		result_out2414<=result2414;
		result_out2415<=result2415;
		result_out2416<=result2416;
		result_out2417<=result2417;
		result_out2418<=result2418;
		result_out2419<=result2419;
		result_out2420<=result2420;
		result_out2421<=result2421;
		result_out2422<=result2422;
		result_out2423<=result2423;
		result_out2424<=result2424;
		result_out2425<=result2425;
		result_out2426<=result2426;
		result_out2427<=result2427;
		result_out2428<=result2428;
		result_out2429<=result2429;
		result_out2430<=result2430;
		result_out2431<=result2431;
		result_out2432<=result2432;
		result_out2433<=result2433;
		result_out2434<=result2434;
		result_out2435<=result2435;
		result_out2436<=result2436;
		result_out2437<=result2437;
		result_out2438<=result2438;
		result_out2439<=result2439;
		result_out2440<=result2440;
		result_out2441<=result2441;
		result_out2442<=result2442;
		result_out2443<=result2443;
		result_out2444<=result2444;
		result_out2445<=result2445;
		result_out2446<=result2446;
		result_out2447<=result2447;
		result_out2448<=result2448;
		result_out2449<=result2449;
		result_out2450<=result2450;
		result_out2451<=result2451;
		result_out2452<=result2452;
		result_out2453<=result2453;
		result_out2454<=result2454;
		result_out2455<=result2455;
		result_out2456<=result2456;
		result_out2457<=result2457;
		result_out2458<=result2458;
		result_out2459<=result2459;
		result_out2460<=result2460;
		result_out2461<=result2461;
		result_out2462<=result2462;
		result_out2463<=result2463;
		result_out2464<=result2464;
		result_out2465<=result2465;
		result_out2466<=result2466;
		result_out2467<=result2467;
		result_out2468<=result2468;
		result_out2469<=result2469;
		result_out2470<=result2470;
		result_out2471<=result2471;
		result_out2472<=result2472;
		result_out2473<=result2473;
		result_out2474<=result2474;
		result_out2475<=result2475;
		result_out2476<=result2476;
		result_out2477<=result2477;
		result_out2478<=result2478;
		result_out2479<=result2479;
		result_out2480<=result2480;
		result_out2481<=result2481;
		result_out2482<=result2482;
		result_out2483<=result2483;
		result_out2484<=result2484;
		result_out2485<=result2485;
		result_out2486<=result2486;
		result_out2487<=result2487;
		result_out2488<=result2488;
		result_out2489<=result2489;
		result_out2490<=result2490;
		result_out2491<=result2491;
		result_out2492<=result2492;
		result_out2493<=result2493;
		result_out2494<=result2494;
		result_out2495<=result2495;
		result_out2496<=result2496;
		result_out2497<=result2497;
		result_out2498<=result2498;
		result_out2499<=result2499;
		result_out2500<=result2500;
		result_out2501<=result2501;
		result_out2502<=result2502;
		result_out2503<=result2503;
		result_out2504<=result2504;
		result_out2505<=result2505;
		result_out2506<=result2506;
		result_out2507<=result2507;
		result_out2508<=result2508;
		result_out2509<=result2509;
		result_out2510<=result2510;
		result_out2511<=result2511;
		result_out2512<=result2512;
		result_out2513<=result2513;
		result_out2514<=result2514;
		result_out2515<=result2515;
		result_out2516<=result2516;
		result_out2517<=result2517;
		result_out2518<=result2518;
		result_out2519<=result2519;
		result_out2520<=result2520;
		result_out2521<=result2521;
		result_out2522<=result2522;
		result_out2523<=result2523;
		result_out2524<=result2524;
		result_out2525<=result2525;
		result_out2526<=result2526;
		result_out2527<=result2527;
		result_out2528<=result2528;
		result_out2529<=result2529;
		result_out2530<=result2530;
		result_out2531<=result2531;
		result_out2532<=result2532;
		result_out2533<=result2533;
		result_out2534<=result2534;
		result_out2535<=result2535;
		result_out2536<=result2536;
		result_out2537<=result2537;
		result_out2538<=result2538;
		result_out2539<=result2539;
		result_out2540<=result2540;
		result_out2541<=result2541;
		result_out2542<=result2542;
		result_out2543<=result2543;
		result_out2544<=result2544;
		result_out2545<=result2545;
		result_out2546<=result2546;
		result_out2547<=result2547;
		result_out2548<=result2548;
		result_out2549<=result2549;
		result_out2550<=result2550;
		result_out2551<=result2551;
		result_out2552<=result2552;
		result_out2553<=result2553;
		result_out2554<=result2554;
		result_out2555<=result2555;
		result_out2556<=result2556;
		result_out2557<=result2557;
		result_out2558<=result2558;
		result_out2559<=result2559;
		result_out2560<=result2560;
		result_out2561<=result2561;
		result_out2562<=result2562;
		result_out2563<=result2563;
		result_out2564<=result2564;
		result_out2565<=result2565;
		result_out2566<=result2566;
		result_out2567<=result2567;
		result_out2568<=result2568;
		result_out2569<=result2569;
		result_out2570<=result2570;
		result_out2571<=result2571;
		result_out2572<=result2572;
		result_out2573<=result2573;
		result_out2574<=result2574;
		result_out2575<=result2575;
		result_out2576<=result2576;
		result_out2577<=result2577;
		result_out2578<=result2578;
		result_out2579<=result2579;
		result_out2580<=result2580;
		result_out2581<=result2581;
		result_out2582<=result2582;
		result_out2583<=result2583;
		result_out2584<=result2584;
		result_out2585<=result2585;
		result_out2586<=result2586;
		result_out2587<=result2587;
		result_out2588<=result2588;
		result_out2589<=result2589;
		result_out2590<=result2590;
		result_out2591<=result2591;
		result_out2592<=result2592;
		result_out2593<=result2593;
		result_out2594<=result2594;
		result_out2595<=result2595;
		result_out2596<=result2596;
		result_out2597<=result2597;
		result_out2598<=result2598;
		result_out2599<=result2599;
		result_out2600<=result2600;
		result_out2601<=result2601;
		result_out2602<=result2602;
		result_out2603<=result2603;
		result_out2604<=result2604;
		result_out2605<=result2605;
		result_out2606<=result2606;
		result_out2607<=result2607;
		result_out2608<=result2608;
		result_out2609<=result2609;
		result_out2610<=result2610;
		result_out2611<=result2611;
		result_out2612<=result2612;
		result_out2613<=result2613;
		result_out2614<=result2614;
		result_out2615<=result2615;
		result_out2616<=result2616;
		result_out2617<=result2617;
		result_out2618<=result2618;
		result_out2619<=result2619;
		result_out2620<=result2620;
		result_out2621<=result2621;
		result_out2622<=result2622;
		result_out2623<=result2623;
		result_out2624<=result2624;
		result_out2625<=result2625;
		result_out2626<=result2626;
		result_out2627<=result2627;
		result_out2628<=result2628;
		result_out2629<=result2629;
		result_out2630<=result2630;
		result_out2631<=result2631;
		result_out2632<=result2632;
		result_out2633<=result2633;
		result_out2634<=result2634;
		result_out2635<=result2635;
		result_out2636<=result2636;
		result_out2637<=result2637;
		result_out2638<=result2638;
		result_out2639<=result2639;
		result_out2640<=result2640;
		result_out2641<=result2641;
		result_out2642<=result2642;
		result_out2643<=result2643;
		result_out2644<=result2644;
		result_out2645<=result2645;
		result_out2646<=result2646;
		result_out2647<=result2647;
		result_out2648<=result2648;
		result_out2649<=result2649;
		result_out2650<=result2650;
		result_out2651<=result2651;
		result_out2652<=result2652;
		result_out2653<=result2653;
		result_out2654<=result2654;
		result_out2655<=result2655;
		result_out2656<=result2656;
		result_out2657<=result2657;
		result_out2658<=result2658;
		result_out2659<=result2659;
		result_out2660<=result2660;
		result_out2661<=result2661;
		result_out2662<=result2662;
		result_out2663<=result2663;
		result_out2664<=result2664;
		result_out2665<=result2665;
		result_out2666<=result2666;
		result_out2667<=result2667;
		result_out2668<=result2668;
		result_out2669<=result2669;
		result_out2670<=result2670;
		result_out2671<=result2671;
		result_out2672<=result2672;
		result_out2673<=result2673;
		result_out2674<=result2674;
		result_out2675<=result2675;
		result_out2676<=result2676;
		result_out2677<=result2677;
		result_out2678<=result2678;
		result_out2679<=result2679;
		result_out2680<=result2680;
		result_out2681<=result2681;
		result_out2682<=result2682;
		result_out2683<=result2683;
		result_out2684<=result2684;
		result_out2685<=result2685;
		result_out2686<=result2686;
		result_out2687<=result2687;
		result_out2688<=result2688;
		result_out2689<=result2689;
		result_out2690<=result2690;
		result_out2691<=result2691;
		result_out2692<=result2692;
		result_out2693<=result2693;
		result_out2694<=result2694;
		result_out2695<=result2695;
		result_out2696<=result2696;
		result_out2697<=result2697;
		result_out2698<=result2698;
		result_out2699<=result2699;
		result_out2700<=result2700;
		result_out2701<=result2701;
		result_out2702<=result2702;
		result_out2703<=result2703;
		result_out2704<=result2704;
		result_out2705<=result2705;
		result_out2706<=result2706;
		result_out2707<=result2707;
		result_out2708<=result2708;
		result_out2709<=result2709;
		result_out2710<=result2710;
		result_out2711<=result2711;
		result_out2712<=result2712;
		result_out2713<=result2713;
		result_out2714<=result2714;
		result_out2715<=result2715;
		result_out2716<=result2716;
		result_out2717<=result2717;
		result_out2718<=result2718;
		result_out2719<=result2719;
		result_out2720<=result2720;
		result_out2721<=result2721;
		result_out2722<=result2722;
		result_out2723<=result2723;
		result_out2724<=result2724;
		result_out2725<=result2725;
		result_out2726<=result2726;
		result_out2727<=result2727;
		result_out2728<=result2728;
		result_out2729<=result2729;
		result_out2730<=result2730;
		result_out2731<=result2731;
		result_out2732<=result2732;
		result_out2733<=result2733;
		result_out2734<=result2734;
		result_out2735<=result2735;
		result_out2736<=result2736;
		result_out2737<=result2737;
		result_out2738<=result2738;
		result_out2739<=result2739;
		result_out2740<=result2740;
		result_out2741<=result2741;
		result_out2742<=result2742;
		result_out2743<=result2743;
		result_out2744<=result2744;
		result_out2745<=result2745;
		result_out2746<=result2746;
		result_out2747<=result2747;
		result_out2748<=result2748;
		result_out2749<=result2749;
		result_out2750<=result2750;
		result_out2751<=result2751;
		result_out2752<=result2752;
		result_out2753<=result2753;
		result_out2754<=result2754;
		result_out2755<=result2755;
		result_out2756<=result2756;
		result_out2757<=result2757;
		result_out2758<=result2758;
		result_out2759<=result2759;
		result_out2760<=result2760;
		result_out2761<=result2761;
		result_out2762<=result2762;
		result_out2763<=result2763;
		result_out2764<=result2764;
		result_out2765<=result2765;
		result_out2766<=result2766;
		result_out2767<=result2767;
		result_out2768<=result2768;
		result_out2769<=result2769;
		result_out2770<=result2770;
		result_out2771<=result2771;
		result_out2772<=result2772;
		result_out2773<=result2773;
		result_out2774<=result2774;
		result_out2775<=result2775;
		result_out2776<=result2776;
		result_out2777<=result2777;
		result_out2778<=result2778;
		result_out2779<=result2779;
		result_out2780<=result2780;
		result_out2781<=result2781;
		result_out2782<=result2782;
		result_out2783<=result2783;
		result_out2784<=result2784;
		result_out2785<=result2785;
		result_out2786<=result2786;
		result_out2787<=result2787;
		result_out2788<=result2788;
		result_out2789<=result2789;
		result_out2790<=result2790;
		result_out2791<=result2791;
		result_out2792<=result2792;
		result_out2793<=result2793;
		result_out2794<=result2794;
		result_out2795<=result2795;
		result_out2796<=result2796;
		result_out2797<=result2797;
		result_out2798<=result2798;
		result_out2799<=result2799;
		result_out2800<=result2800;
		result_out2801<=result2801;
		result_out2802<=result2802;
		result_out2803<=result2803;
		result_out2804<=result2804;
		result_out2805<=result2805;
		result_out2806<=result2806;
		result_out2807<=result2807;
		result_out2808<=result2808;
		result_out2809<=result2809;
		result_out2810<=result2810;
		result_out2811<=result2811;
		result_out2812<=result2812;
		result_out2813<=result2813;
		result_out2814<=result2814;
		result_out2815<=result2815;
		result_out2816<=result2816;
		result_out2817<=result2817;
		result_out2818<=result2818;
		result_out2819<=result2819;
		result_out2820<=result2820;
		result_out2821<=result2821;
		result_out2822<=result2822;
		result_out2823<=result2823;
		result_out2824<=result2824;
		result_out2825<=result2825;
		result_out2826<=result2826;
		result_out2827<=result2827;
		result_out2828<=result2828;
		result_out2829<=result2829;
		result_out2830<=result2830;
		result_out2831<=result2831;
		result_out2832<=result2832;
		result_out2833<=result2833;
		result_out2834<=result2834;
		result_out2835<=result2835;
		result_out2836<=result2836;
		result_out2837<=result2837;
		result_out2838<=result2838;
		result_out2839<=result2839;
		result_out2840<=result2840;
		result_out2841<=result2841;
		result_out2842<=result2842;
		result_out2843<=result2843;
		result_out2844<=result2844;
		result_out2845<=result2845;
		result_out2846<=result2846;
		result_out2847<=result2847;
		result_out2848<=result2848;
		result_out2849<=result2849;
		result_out2850<=result2850;
		result_out2851<=result2851;
		result_out2852<=result2852;
		result_out2853<=result2853;
		result_out2854<=result2854;
		result_out2855<=result2855;
		result_out2856<=result2856;
		result_out2857<=result2857;
		result_out2858<=result2858;
		result_out2859<=result2859;
		result_out2860<=result2860;
		result_out2861<=result2861;
		result_out2862<=result2862;
		result_out2863<=result2863;
		result_out2864<=result2864;
		result_out2865<=result2865;
		result_out2866<=result2866;
		result_out2867<=result2867;
		result_out2868<=result2868;
		result_out2869<=result2869;
		result_out2870<=result2870;
		result_out2871<=result2871;
		result_out2872<=result2872;
		result_out2873<=result2873;
		result_out2874<=result2874;
		result_out2875<=result2875;
		result_out2876<=result2876;
		result_out2877<=result2877;
		result_out2878<=result2878;
		result_out2879<=result2879;
		result_out2880<=result2880;
		result_out2881<=result2881;
		result_out2882<=result2882;
		result_out2883<=result2883;
		result_out2884<=result2884;
		result_out2885<=result2885;
		result_out2886<=result2886;
		result_out2887<=result2887;
		result_out2888<=result2888;
		result_out2889<=result2889;
		result_out2890<=result2890;
		result_out2891<=result2891;
		result_out2892<=result2892;
		result_out2893<=result2893;
		result_out2894<=result2894;
		result_out2895<=result2895;
		result_out2896<=result2896;
		result_out2897<=result2897;
		result_out2898<=result2898;
		result_out2899<=result2899;
		result_out2900<=result2900;
		result_out2901<=result2901;
		result_out2902<=result2902;
		result_out2903<=result2903;
		result_out2904<=result2904;
		result_out2905<=result2905;
		result_out2906<=result2906;
		result_out2907<=result2907;
		result_out2908<=result2908;
		result_out2909<=result2909;
		result_out2910<=result2910;
		result_out2911<=result2911;
		result_out2912<=result2912;
		result_out2913<=result2913;
		result_out2914<=result2914;
		result_out2915<=result2915;
		result_out2916<=result2916;
		result_out2917<=result2917;
		result_out2918<=result2918;
		result_out2919<=result2919;
		result_out2920<=result2920;
		result_out2921<=result2921;
		result_out2922<=result2922;
		result_out2923<=result2923;
		result_out2924<=result2924;
		result_out2925<=result2925;
		result_out2926<=result2926;
		result_out2927<=result2927;
		result_out2928<=result2928;
		result_out2929<=result2929;
		result_out2930<=result2930;
		result_out2931<=result2931;
		result_out2932<=result2932;
		result_out2933<=result2933;
		result_out2934<=result2934;
		result_out2935<=result2935;
		result_out2936<=result2936;
		result_out2937<=result2937;
		result_out2938<=result2938;
		result_out2939<=result2939;
		result_out2940<=result2940;
		result_out2941<=result2941;
		result_out2942<=result2942;
		result_out2943<=result2943;
		result_out2944<=result2944;
		result_out2945<=result2945;
		result_out2946<=result2946;
		result_out2947<=result2947;
		result_out2948<=result2948;
		result_out2949<=result2949;
		result_out2950<=result2950;
		result_out2951<=result2951;
		result_out2952<=result2952;
		result_out2953<=result2953;
		result_out2954<=result2954;
		result_out2955<=result2955;
		result_out2956<=result2956;
		result_out2957<=result2957;
		result_out2958<=result2958;
		result_out2959<=result2959;
		result_out2960<=result2960;
		result_out2961<=result2961;
		result_out2962<=result2962;
		result_out2963<=result2963;
		result_out2964<=result2964;
		result_out2965<=result2965;
		result_out2966<=result2966;
		result_out2967<=result2967;
		result_out2968<=result2968;
		result_out2969<=result2969;
		result_out2970<=result2970;
		result_out2971<=result2971;
		result_out2972<=result2972;
		result_out2973<=result2973;
		result_out2974<=result2974;
		result_out2975<=result2975;
		result_out2976<=result2976;
		result_out2977<=result2977;
		result_out2978<=result2978;
		result_out2979<=result2979;
		result_out2980<=result2980;
		result_out2981<=result2981;
		result_out2982<=result2982;
		result_out2983<=result2983;
		result_out2984<=result2984;
		result_out2985<=result2985;
		result_out2986<=result2986;
		result_out2987<=result2987;
		result_out2988<=result2988;
		result_out2989<=result2989;
		result_out2990<=result2990;
		result_out2991<=result2991;
		result_out2992<=result2992;
		result_out2993<=result2993;
		result_out2994<=result2994;
		result_out2995<=result2995;
		result_out2996<=result2996;
		result_out2997<=result2997;
		result_out2998<=result2998;
		result_out2999<=result2999;
		result_out3000<=result3000;
		result_out3001<=result3001;
		result_out3002<=result3002;
		result_out3003<=result3003;
		result_out3004<=result3004;
		result_out3005<=result3005;
		result_out3006<=result3006;
		result_out3007<=result3007;
		result_out3008<=result3008;
		result_out3009<=result3009;
		result_out3010<=result3010;
		result_out3011<=result3011;
		result_out3012<=result3012;
		result_out3013<=result3013;
		result_out3014<=result3014;
		result_out3015<=result3015;
		result_out3016<=result3016;
		result_out3017<=result3017;
		result_out3018<=result3018;
		result_out3019<=result3019;
		result_out3020<=result3020;
		result_out3021<=result3021;
		result_out3022<=result3022;
		result_out3023<=result3023;
		result_out3024<=result3024;
		result_out3025<=result3025;
		result_out3026<=result3026;
		result_out3027<=result3027;
		result_out3028<=result3028;
		result_out3029<=result3029;
		result_out3030<=result3030;
		result_out3031<=result3031;
		result_out3032<=result3032;
		result_out3033<=result3033;
		result_out3034<=result3034;
		result_out3035<=result3035;
		result_out3036<=result3036;
		result_out3037<=result3037;
		result_out3038<=result3038;
		result_out3039<=result3039;
		result_out3040<=result3040;
		result_out3041<=result3041;
		result_out3042<=result3042;
		result_out3043<=result3043;
		result_out3044<=result3044;
		result_out3045<=result3045;
		result_out3046<=result3046;
		result_out3047<=result3047;
		result_out3048<=result3048;
		result_out3049<=result3049;
		result_out3050<=result3050;
		result_out3051<=result3051;
		result_out3052<=result3052;
		result_out3053<=result3053;
		result_out3054<=result3054;
		result_out3055<=result3055;
		result_out3056<=result3056;
		result_out3057<=result3057;
		result_out3058<=result3058;
		result_out3059<=result3059;
		result_out3060<=result3060;
		result_out3061<=result3061;
		result_out3062<=result3062;
		result_out3063<=result3063;
		result_out3064<=result3064;
		result_out3065<=result3065;
		result_out3066<=result3066;
		result_out3067<=result3067;
		result_out3068<=result3068;
		result_out3069<=result3069;
		result_out3070<=result3070;
		result_out3071<=result3071;
		result_out3072<=result3072;
		result_out3073<=result3073;
		result_out3074<=result3074;
		result_out3075<=result3075;
		result_out3076<=result3076;
		result_out3077<=result3077;
		result_out3078<=result3078;
		result_out3079<=result3079;
		result_out3080<=result3080;
		result_out3081<=result3081;
		result_out3082<=result3082;
		result_out3083<=result3083;
		result_out3084<=result3084;
		result_out3085<=result3085;
		result_out3086<=result3086;
		result_out3087<=result3087;
		result_out3088<=result3088;
		result_out3089<=result3089;
		result_out3090<=result3090;
		result_out3091<=result3091;
		result_out3092<=result3092;
		result_out3093<=result3093;
		result_out3094<=result3094;
		result_out3095<=result3095;
		result_out3096<=result3096;
		result_out3097<=result3097;
		result_out3098<=result3098;
		result_out3099<=result3099;
		result_out3100<=result3100;
		result_out3101<=result3101;
		result_out3102<=result3102;
		result_out3103<=result3103;
		result_out3104<=result3104;
		result_out3105<=result3105;
		result_out3106<=result3106;
		result_out3107<=result3107;
		result_out3108<=result3108;
		result_out3109<=result3109;
		result_out3110<=result3110;
		result_out3111<=result3111;
		result_out3112<=result3112;
		result_out3113<=result3113;
		result_out3114<=result3114;
		result_out3115<=result3115;
		result_out3116<=result3116;
		result_out3117<=result3117;
		result_out3118<=result3118;
		result_out3119<=result3119;
		result_out3120<=result3120;
		result_out3121<=result3121;
		result_out3122<=result3122;
		result_out3123<=result3123;
		result_out3124<=result3124;
		result_out3125<=result3125;
		result_out3126<=result3126;
		result_out3127<=result3127;
		result_out3128<=result3128;
		result_out3129<=result3129;
		result_out3130<=result3130;
		result_out3131<=result3131;
		result_out3132<=result3132;
		result_out3133<=result3133;
		result_out3134<=result3134;
		result_out3135<=result3135;
		result_out3136<=result3136;
		result_out3137<=result3137;
		result_out3138<=result3138;
		result_out3139<=result3139;
		result_out3140<=result3140;
		result_out3141<=result3141;
		result_out3142<=result3142;
		result_out3143<=result3143;
		result_out3144<=result3144;
		result_out3145<=result3145;
		result_out3146<=result3146;
		result_out3147<=result3147;
		result_out3148<=result3148;
		result_out3149<=result3149;
		result_out3150<=result3150;
		result_out3151<=result3151;
		result_out3152<=result3152;
		result_out3153<=result3153;
		result_out3154<=result3154;
		result_out3155<=result3155;
		result_out3156<=result3156;
		result_out3157<=result3157;
		result_out3158<=result3158;
		result_out3159<=result3159;
		result_out3160<=result3160;
		result_out3161<=result3161;
		result_out3162<=result3162;
		result_out3163<=result3163;
		result_out3164<=result3164;
		result_out3165<=result3165;
		result_out3166<=result3166;
		result_out3167<=result3167;
		result_out3168<=result3168;
		result_out3169<=result3169;
		result_out3170<=result3170;
		result_out3171<=result3171;
		result_out3172<=result3172;
		result_out3173<=result3173;
		result_out3174<=result3174;
		result_out3175<=result3175;
		result_out3176<=result3176;
		result_out3177<=result3177;
		result_out3178<=result3178;
		result_out3179<=result3179;
		result_out3180<=result3180;
		result_out3181<=result3181;
		result_out3182<=result3182;
		result_out3183<=result3183;
		result_out3184<=result3184;
		result_out3185<=result3185;
		result_out3186<=result3186;
		result_out3187<=result3187;
		result_out3188<=result3188;
		result_out3189<=result3189;
		result_out3190<=result3190;
		result_out3191<=result3191;
		result_out3192<=result3192;
		result_out3193<=result3193;
		result_out3194<=result3194;
		result_out3195<=result3195;
		result_out3196<=result3196;
		result_out3197<=result3197;
		result_out3198<=result3198;
		result_out3199<=result3199;
		result_out3200<=result3200;
		result_out3201<=result3201;
		result_out3202<=result3202;
		result_out3203<=result3203;
		result_out3204<=result3204;
		result_out3205<=result3205;
		result_out3206<=result3206;
		result_out3207<=result3207;
		result_out3208<=result3208;
		result_out3209<=result3209;
		result_out3210<=result3210;
		result_out3211<=result3211;
		result_out3212<=result3212;
		result_out3213<=result3213;
		result_out3214<=result3214;
		result_out3215<=result3215;
		result_out3216<=result3216;
		result_out3217<=result3217;
		result_out3218<=result3218;
		result_out3219<=result3219;
		result_out3220<=result3220;
		result_out3221<=result3221;
		result_out3222<=result3222;
		result_out3223<=result3223;
		result_out3224<=result3224;
		result_out3225<=result3225;
		result_out3226<=result3226;
		result_out3227<=result3227;
		result_out3228<=result3228;
		result_out3229<=result3229;
		result_out3230<=result3230;
		result_out3231<=result3231;
		result_out3232<=result3232;
		result_out3233<=result3233;
		result_out3234<=result3234;
		result_out3235<=result3235;
		result_out3236<=result3236;
		result_out3237<=result3237;
		result_out3238<=result3238;
		result_out3239<=result3239;
		result_out3240<=result3240;
		result_out3241<=result3241;
		result_out3242<=result3242;
		result_out3243<=result3243;
		result_out3244<=result3244;
		result_out3245<=result3245;
		result_out3246<=result3246;
		result_out3247<=result3247;
		result_out3248<=result3248;
		result_out3249<=result3249;
		result_out3250<=result3250;
		result_out3251<=result3251;
		result_out3252<=result3252;
		result_out3253<=result3253;
		result_out3254<=result3254;
		result_out3255<=result3255;
		result_out3256<=result3256;
		result_out3257<=result3257;
		result_out3258<=result3258;
		result_out3259<=result3259;
		result_out3260<=result3260;
		result_out3261<=result3261;
		result_out3262<=result3262;
		result_out3263<=result3263;
		result_out3264<=result3264;
		result_out3265<=result3265;
		result_out3266<=result3266;
		result_out3267<=result3267;
		result_out3268<=result3268;
		result_out3269<=result3269;
		result_out3270<=result3270;
		result_out3271<=result3271;
		result_out3272<=result3272;
		result_out3273<=result3273;
		result_out3274<=result3274;
		result_out3275<=result3275;
		result_out3276<=result3276;
		result_out3277<=result3277;
		result_out3278<=result3278;
		result_out3279<=result3279;
		result_out3280<=result3280;
		result_out3281<=result3281;
		result_out3282<=result3282;
		result_out3283<=result3283;
		result_out3284<=result3284;
		result_out3285<=result3285;
		result_out3286<=result3286;
		result_out3287<=result3287;
		result_out3288<=result3288;
		result_out3289<=result3289;
		result_out3290<=result3290;
		result_out3291<=result3291;
		result_out3292<=result3292;
		result_out3293<=result3293;
		result_out3294<=result3294;
		result_out3295<=result3295;
		result_out3296<=result3296;
		result_out3297<=result3297;
		result_out3298<=result3298;
		result_out3299<=result3299;
		result_out3300<=result3300;
		result_out3301<=result3301;
		result_out3302<=result3302;
		result_out3303<=result3303;
		result_out3304<=result3304;
		result_out3305<=result3305;
		result_out3306<=result3306;
		result_out3307<=result3307;
		result_out3308<=result3308;
		result_out3309<=result3309;
		result_out3310<=result3310;
		result_out3311<=result3311;
		result_out3312<=result3312;
		result_out3313<=result3313;
		result_out3314<=result3314;
		result_out3315<=result3315;
		result_out3316<=result3316;
		result_out3317<=result3317;
		result_out3318<=result3318;
		result_out3319<=result3319;
		result_out3320<=result3320;
		result_out3321<=result3321;
		result_out3322<=result3322;
		result_out3323<=result3323;
		result_out3324<=result3324;
		result_out3325<=result3325;
		result_out3326<=result3326;
		result_out3327<=result3327;
		result_out3328<=result3328;
		result_out3329<=result3329;
		result_out3330<=result3330;
		result_out3331<=result3331;
		result_out3332<=result3332;
		result_out3333<=result3333;
		result_out3334<=result3334;
		result_out3335<=result3335;
		result_out3336<=result3336;
		result_out3337<=result3337;
		result_out3338<=result3338;
		result_out3339<=result3339;
		result_out3340<=result3340;
		result_out3341<=result3341;
		result_out3342<=result3342;
		result_out3343<=result3343;
		result_out3344<=result3344;
		result_out3345<=result3345;
		result_out3346<=result3346;
		result_out3347<=result3347;
		result_out3348<=result3348;
		result_out3349<=result3349;
		result_out3350<=result3350;
		result_out3351<=result3351;
		result_out3352<=result3352;
		result_out3353<=result3353;
		result_out3354<=result3354;
		result_out3355<=result3355;
		result_out3356<=result3356;
		result_out3357<=result3357;
		result_out3358<=result3358;
		result_out3359<=result3359;
		result_out3360<=result3360;
		result_out3361<=result3361;
		result_out3362<=result3362;
		result_out3363<=result3363;
		result_out3364<=result3364;
		result_out3365<=result3365;
		result_out3366<=result3366;
		result_out3367<=result3367;
		result_out3368<=result3368;
		result_out3369<=result3369;
		result_out3370<=result3370;
		result_out3371<=result3371;
		result_out3372<=result3372;
		result_out3373<=result3373;
		result_out3374<=result3374;
		result_out3375<=result3375;
		result_out3376<=result3376;
		result_out3377<=result3377;
		result_out3378<=result3378;
		result_out3379<=result3379;
		result_out3380<=result3380;
		result_out3381<=result3381;
		result_out3382<=result3382;
		result_out3383<=result3383;
		result_out3384<=result3384;
		result_out3385<=result3385;
		result_out3386<=result3386;
		result_out3387<=result3387;
		result_out3388<=result3388;
		result_out3389<=result3389;
		result_out3390<=result3390;
		result_out3391<=result3391;
		result_out3392<=result3392;
		result_out3393<=result3393;
		result_out3394<=result3394;
		result_out3395<=result3395;
		result_out3396<=result3396;
		result_out3397<=result3397;
		result_out3398<=result3398;
		result_out3399<=result3399;
		result_out3400<=result3400;
		result_out3401<=result3401;
		result_out3402<=result3402;
		result_out3403<=result3403;
		result_out3404<=result3404;
		result_out3405<=result3405;
		result_out3406<=result3406;
		result_out3407<=result3407;
		result_out3408<=result3408;
		result_out3409<=result3409;
		result_out3410<=result3410;
		result_out3411<=result3411;
		result_out3412<=result3412;
		result_out3413<=result3413;
		result_out3414<=result3414;
		result_out3415<=result3415;
		result_out3416<=result3416;
		result_out3417<=result3417;
		result_out3418<=result3418;
		result_out3419<=result3419;
		result_out3420<=result3420;
		result_out3421<=result3421;
		result_out3422<=result3422;
		result_out3423<=result3423;
		result_out3424<=result3424;
		result_out3425<=result3425;
		result_out3426<=result3426;
		result_out3427<=result3427;
		result_out3428<=result3428;
		result_out3429<=result3429;
		result_out3430<=result3430;
		result_out3431<=result3431;
		result_out3432<=result3432;
		result_out3433<=result3433;
		result_out3434<=result3434;
		result_out3435<=result3435;
		result_out3436<=result3436;
		result_out3437<=result3437;
		result_out3438<=result3438;
		result_out3439<=result3439;
		result_out3440<=result3440;
		result_out3441<=result3441;
		result_out3442<=result3442;
		result_out3443<=result3443;
		result_out3444<=result3444;
		result_out3445<=result3445;
		result_out3446<=result3446;
		result_out3447<=result3447;
		result_out3448<=result3448;
		result_out3449<=result3449;
		result_out3450<=result3450;
		result_out3451<=result3451;
		result_out3452<=result3452;
		result_out3453<=result3453;
		result_out3454<=result3454;
		result_out3455<=result3455;
		result_out3456<=result3456;
		result_out3457<=result3457;
		result_out3458<=result3458;
		result_out3459<=result3459;
		result_out3460<=result3460;
		result_out3461<=result3461;
		result_out3462<=result3462;
		result_out3463<=result3463;
		result_out3464<=result3464;
		result_out3465<=result3465;
		result_out3466<=result3466;
		result_out3467<=result3467;
		result_out3468<=result3468;
		result_out3469<=result3469;
		result_out3470<=result3470;
		result_out3471<=result3471;
		result_out3472<=result3472;
		result_out3473<=result3473;
		result_out3474<=result3474;
		result_out3475<=result3475;
		result_out3476<=result3476;
		result_out3477<=result3477;
		result_out3478<=result3478;
		result_out3479<=result3479;
		result_out3480<=result3480;
		result_out3481<=result3481;
		result_out3482<=result3482;
		result_out3483<=result3483;
		result_out3484<=result3484;
		result_out3485<=result3485;
		result_out3486<=result3486;
		result_out3487<=result3487;
		result_out3488<=result3488;
		result_out3489<=result3489;
		result_out3490<=result3490;
		result_out3491<=result3491;
		result_out3492<=result3492;
		result_out3493<=result3493;
		result_out3494<=result3494;
		result_out3495<=result3495;
		result_out3496<=result3496;
		result_out3497<=result3497;
		result_out3498<=result3498;
		result_out3499<=result3499;
		result_out3500<=result3500;
		result_out3501<=result3501;
		result_out3502<=result3502;
		result_out3503<=result3503;
		result_out3504<=result3504;
		result_out3505<=result3505;
		result_out3506<=result3506;
		result_out3507<=result3507;
		result_out3508<=result3508;
		result_out3509<=result3509;
		result_out3510<=result3510;
		result_out3511<=result3511;
		result_out3512<=result3512;
		result_out3513<=result3513;
		result_out3514<=result3514;
		result_out3515<=result3515;
		result_out3516<=result3516;
		result_out3517<=result3517;
		result_out3518<=result3518;
		result_out3519<=result3519;
		result_out3520<=result3520;
		result_out3521<=result3521;
		result_out3522<=result3522;
		result_out3523<=result3523;
		result_out3524<=result3524;
		result_out3525<=result3525;
		result_out3526<=result3526;
		result_out3527<=result3527;
		result_out3528<=result3528;
		result_out3529<=result3529;
		result_out3530<=result3530;
		result_out3531<=result3531;
		result_out3532<=result3532;
		result_out3533<=result3533;
		result_out3534<=result3534;
		result_out3535<=result3535;
		result_out3536<=result3536;
		result_out3537<=result3537;
		result_out3538<=result3538;
		result_out3539<=result3539;
		result_out3540<=result3540;
		result_out3541<=result3541;
		result_out3542<=result3542;
		result_out3543<=result3543;
		result_out3544<=result3544;
		result_out3545<=result3545;
		result_out3546<=result3546;
		result_out3547<=result3547;
		result_out3548<=result3548;
		result_out3549<=result3549;
		result_out3550<=result3550;
		result_out3551<=result3551;
		result_out3552<=result3552;
		result_out3553<=result3553;
		result_out3554<=result3554;
		result_out3555<=result3555;
		result_out3556<=result3556;
		result_out3557<=result3557;
		result_out3558<=result3558;
		result_out3559<=result3559;
		result_out3560<=result3560;
		result_out3561<=result3561;
		result_out3562<=result3562;
		result_out3563<=result3563;
		result_out3564<=result3564;
		result_out3565<=result3565;
		result_out3566<=result3566;
		result_out3567<=result3567;
		result_out3568<=result3568;
		result_out3569<=result3569;
		result_out3570<=result3570;
		result_out3571<=result3571;
		result_out3572<=result3572;
		result_out3573<=result3573;
		result_out3574<=result3574;
		result_out3575<=result3575;
		result_out3576<=result3576;
		result_out3577<=result3577;
		result_out3578<=result3578;
		result_out3579<=result3579;
		result_out3580<=result3580;
		result_out3581<=result3581;
		result_out3582<=result3582;
		result_out3583<=result3583;
		result_out3584<=result3584;
		result_out3585<=result3585;
		result_out3586<=result3586;
		result_out3587<=result3587;
		result_out3588<=result3588;
		result_out3589<=result3589;
		result_out3590<=result3590;
		result_out3591<=result3591;
		result_out3592<=result3592;
		result_out3593<=result3593;
		result_out3594<=result3594;
		result_out3595<=result3595;
		result_out3596<=result3596;
		result_out3597<=result3597;
		result_out3598<=result3598;
		result_out3599<=result3599;
		result_out3600<=result3600;
		result_out3601<=result3601;
		result_out3602<=result3602;
		result_out3603<=result3603;
		result_out3604<=result3604;
		result_out3605<=result3605;
		result_out3606<=result3606;
		result_out3607<=result3607;
		result_out3608<=result3608;
		result_out3609<=result3609;
		result_out3610<=result3610;
		result_out3611<=result3611;
		result_out3612<=result3612;
		result_out3613<=result3613;
		result_out3614<=result3614;
		result_out3615<=result3615;
		result_out3616<=result3616;
		result_out3617<=result3617;
		result_out3618<=result3618;
		result_out3619<=result3619;
		result_out3620<=result3620;
		result_out3621<=result3621;
		result_out3622<=result3622;
		result_out3623<=result3623;
		result_out3624<=result3624;
		result_out3625<=result3625;
		result_out3626<=result3626;
		result_out3627<=result3627;
		result_out3628<=result3628;
		result_out3629<=result3629;
		result_out3630<=result3630;
		result_out3631<=result3631;
		result_out3632<=result3632;
		result_out3633<=result3633;
		result_out3634<=result3634;
		result_out3635<=result3635;
		result_out3636<=result3636;
		result_out3637<=result3637;
		result_out3638<=result3638;
		result_out3639<=result3639;
		result_out3640<=result3640;
		result_out3641<=result3641;
		result_out3642<=result3642;
		result_out3643<=result3643;
		result_out3644<=result3644;
		result_out3645<=result3645;
		result_out3646<=result3646;
		result_out3647<=result3647;
		result_out3648<=result3648;
		result_out3649<=result3649;
		result_out3650<=result3650;
		result_out3651<=result3651;
		result_out3652<=result3652;
		result_out3653<=result3653;
		result_out3654<=result3654;
		result_out3655<=result3655;
		result_out3656<=result3656;
		result_out3657<=result3657;
		result_out3658<=result3658;
		result_out3659<=result3659;
		result_out3660<=result3660;
		result_out3661<=result3661;
		result_out3662<=result3662;
		result_out3663<=result3663;
		result_out3664<=result3664;
		result_out3665<=result3665;
		result_out3666<=result3666;
		result_out3667<=result3667;
		result_out3668<=result3668;
		result_out3669<=result3669;
		result_out3670<=result3670;
		result_out3671<=result3671;
		result_out3672<=result3672;
		result_out3673<=result3673;
		result_out3674<=result3674;
		result_out3675<=result3675;
		result_out3676<=result3676;
		result_out3677<=result3677;
		result_out3678<=result3678;
		result_out3679<=result3679;
		result_out3680<=result3680;
		result_out3681<=result3681;
		result_out3682<=result3682;
		result_out3683<=result3683;
		result_out3684<=result3684;
		result_out3685<=result3685;
		result_out3686<=result3686;
		result_out3687<=result3687;
		result_out3688<=result3688;
		result_out3689<=result3689;
		result_out3690<=result3690;
		result_out3691<=result3691;
		result_out3692<=result3692;
		result_out3693<=result3693;
		result_out3694<=result3694;
		result_out3695<=result3695;
		result_out3696<=result3696;
		result_out3697<=result3697;
		result_out3698<=result3698;
		result_out3699<=result3699;
		result_out3700<=result3700;
		result_out3701<=result3701;
		result_out3702<=result3702;
		result_out3703<=result3703;
		result_out3704<=result3704;
		result_out3705<=result3705;
		result_out3706<=result3706;
		result_out3707<=result3707;
		result_out3708<=result3708;
		result_out3709<=result3709;
		result_out3710<=result3710;
		result_out3711<=result3711;
		result_out3712<=result3712;
		result_out3713<=result3713;
		result_out3714<=result3714;
		result_out3715<=result3715;
		result_out3716<=result3716;
		result_out3717<=result3717;
		result_out3718<=result3718;
		result_out3719<=result3719;
		result_out3720<=result3720;
		result_out3721<=result3721;
		result_out3722<=result3722;
		result_out3723<=result3723;
		result_out3724<=result3724;
		result_out3725<=result3725;
		result_out3726<=result3726;
		result_out3727<=result3727;
		result_out3728<=result3728;
		result_out3729<=result3729;
		result_out3730<=result3730;
		result_out3731<=result3731;
		result_out3732<=result3732;
		result_out3733<=result3733;
		result_out3734<=result3734;
		result_out3735<=result3735;
		result_out3736<=result3736;
		result_out3737<=result3737;
		result_out3738<=result3738;
		result_out3739<=result3739;
		result_out3740<=result3740;
		result_out3741<=result3741;
		result_out3742<=result3742;
		result_out3743<=result3743;
		result_out3744<=result3744;
		result_out3745<=result3745;
		result_out3746<=result3746;
		result_out3747<=result3747;
		result_out3748<=result3748;
		result_out3749<=result3749;
		result_out3750<=result3750;
		result_out3751<=result3751;
		result_out3752<=result3752;
		result_out3753<=result3753;
		result_out3754<=result3754;
		result_out3755<=result3755;
		result_out3756<=result3756;
		result_out3757<=result3757;
		result_out3758<=result3758;
		result_out3759<=result3759;
		result_out3760<=result3760;
		result_out3761<=result3761;
		result_out3762<=result3762;
		result_out3763<=result3763;
		result_out3764<=result3764;
		result_out3765<=result3765;
		result_out3766<=result3766;
		result_out3767<=result3767;
		result_out3768<=result3768;
		result_out3769<=result3769;
		result_out3770<=result3770;
		result_out3771<=result3771;
		result_out3772<=result3772;
		result_out3773<=result3773;
		result_out3774<=result3774;
		result_out3775<=result3775;
		result_out3776<=result3776;
		result_out3777<=result3777;
		result_out3778<=result3778;
		result_out3779<=result3779;
		result_out3780<=result3780;
		result_out3781<=result3781;
		result_out3782<=result3782;
		result_out3783<=result3783;
		result_out3784<=result3784;
		result_out3785<=result3785;
		result_out3786<=result3786;
		result_out3787<=result3787;
		result_out3788<=result3788;
		result_out3789<=result3789;
		result_out3790<=result3790;
		result_out3791<=result3791;
		result_out3792<=result3792;
		result_out3793<=result3793;
		result_out3794<=result3794;
		result_out3795<=result3795;
		result_out3796<=result3796;
		result_out3797<=result3797;
		result_out3798<=result3798;
		result_out3799<=result3799;
		result_out3800<=result3800;
		result_out3801<=result3801;
		result_out3802<=result3802;
		result_out3803<=result3803;
		result_out3804<=result3804;
		result_out3805<=result3805;
		result_out3806<=result3806;
		result_out3807<=result3807;
		result_out3808<=result3808;
		result_out3809<=result3809;
		result_out3810<=result3810;
		result_out3811<=result3811;
		result_out3812<=result3812;
		result_out3813<=result3813;
		result_out3814<=result3814;
		result_out3815<=result3815;
		result_out3816<=result3816;
		result_out3817<=result3817;
		result_out3818<=result3818;
		result_out3819<=result3819;
		result_out3820<=result3820;
		result_out3821<=result3821;
		result_out3822<=result3822;
		result_out3823<=result3823;
		result_out3824<=result3824;
		result_out3825<=result3825;
		result_out3826<=result3826;
		result_out3827<=result3827;
		result_out3828<=result3828;
		result_out3829<=result3829;
		result_out3830<=result3830;
		result_out3831<=result3831;
		result_out3832<=result3832;
		result_out3833<=result3833;
		result_out3834<=result3834;
		result_out3835<=result3835;
		result_out3836<=result3836;
		result_out3837<=result3837;
		result_out3838<=result3838;
		result_out3839<=result3839;
		result_out3840<=result3840;
		result_out3841<=result3841;
		result_out3842<=result3842;
		result_out3843<=result3843;
		result_out3844<=result3844;
		result_out3845<=result3845;
		result_out3846<=result3846;
		result_out3847<=result3847;
		result_out3848<=result3848;
		result_out3849<=result3849;
		result_out3850<=result3850;
		result_out3851<=result3851;
		result_out3852<=result3852;
		result_out3853<=result3853;
		result_out3854<=result3854;
		result_out3855<=result3855;
		result_out3856<=result3856;
		result_out3857<=result3857;
		result_out3858<=result3858;
		result_out3859<=result3859;
		result_out3860<=result3860;
		result_out3861<=result3861;
		result_out3862<=result3862;
		result_out3863<=result3863;
		result_out3864<=result3864;
		result_out3865<=result3865;
		result_out3866<=result3866;
		result_out3867<=result3867;
		result_out3868<=result3868;
		result_out3869<=result3869;
		result_out3870<=result3870;
		result_out3871<=result3871;
		result_out3872<=result3872;
		result_out3873<=result3873;
		result_out3874<=result3874;
		result_out3875<=result3875;
		result_out3876<=result3876;
		result_out3877<=result3877;
		result_out3878<=result3878;
		result_out3879<=result3879;
		result_out3880<=result3880;
		result_out3881<=result3881;
		result_out3882<=result3882;
		result_out3883<=result3883;
		result_out3884<=result3884;
		result_out3885<=result3885;
		result_out3886<=result3886;
		result_out3887<=result3887;
		result_out3888<=result3888;
		result_out3889<=result3889;
		result_out3890<=result3890;
		result_out3891<=result3891;
		result_out3892<=result3892;
		result_out3893<=result3893;
		result_out3894<=result3894;
		result_out3895<=result3895;
		result_out3896<=result3896;
		result_out3897<=result3897;
		result_out3898<=result3898;
		result_out3899<=result3899;
		result_out3900<=result3900;
		result_out3901<=result3901;
		result_out3902<=result3902;
		result_out3903<=result3903;
		result_out3904<=result3904;
		result_out3905<=result3905;
		result_out3906<=result3906;
		result_out3907<=result3907;
		result_out3908<=result3908;
		result_out3909<=result3909;
		result_out3910<=result3910;
		result_out3911<=result3911;
		result_out3912<=result3912;
		result_out3913<=result3913;
		result_out3914<=result3914;
		result_out3915<=result3915;
		result_out3916<=result3916;
		result_out3917<=result3917;
		result_out3918<=result3918;
		result_out3919<=result3919;
		result_out3920<=result3920;
		result_out3921<=result3921;
		result_out3922<=result3922;
		result_out3923<=result3923;
		result_out3924<=result3924;
		result_out3925<=result3925;
		result_out3926<=result3926;
		result_out3927<=result3927;
		result_out3928<=result3928;
		result_out3929<=result3929;
		result_out3930<=result3930;
		result_out3931<=result3931;
		result_out3932<=result3932;
		result_out3933<=result3933;
		result_out3934<=result3934;
		result_out3935<=result3935;
		result_out3936<=result3936;
		result_out3937<=result3937;
		result_out3938<=result3938;
		result_out3939<=result3939;
		result_out3940<=result3940;
		result_out3941<=result3941;
		result_out3942<=result3942;
		result_out3943<=result3943;
		result_out3944<=result3944;
		result_out3945<=result3945;
		result_out3946<=result3946;
		result_out3947<=result3947;
		result_out3948<=result3948;
		result_out3949<=result3949;
		result_out3950<=result3950;
		result_out3951<=result3951;
		result_out3952<=result3952;
		result_out3953<=result3953;
		result_out3954<=result3954;
		result_out3955<=result3955;
		result_out3956<=result3956;
		result_out3957<=result3957;
		result_out3958<=result3958;
		result_out3959<=result3959;
		result_out3960<=result3960;
		result_out3961<=result3961;
		result_out3962<=result3962;
		result_out3963<=result3963;
		result_out3964<=result3964;
		result_out3965<=result3965;
		result_out3966<=result3966;
		result_out3967<=result3967;
		result_out3968<=result3968;
		result_out3969<=result3969;
		result_out3970<=result3970;
		result_out3971<=result3971;
		result_out3972<=result3972;
		result_out3973<=result3973;
		result_out3974<=result3974;
		result_out3975<=result3975;
		result_out3976<=result3976;
		result_out3977<=result3977;
		result_out3978<=result3978;
		result_out3979<=result3979;
		result_out3980<=result3980;
		result_out3981<=result3981;
		result_out3982<=result3982;
		result_out3983<=result3983;
		result_out3984<=result3984;
		result_out3985<=result3985;
		result_out3986<=result3986;
		result_out3987<=result3987;
		result_out3988<=result3988;
		result_out3989<=result3989;
		result_out3990<=result3990;
		result_out3991<=result3991;
		result_out3992<=result3992;
		result_out3993<=result3993;
		result_out3994<=result3994;
		result_out3995<=result3995;
		result_out3996<=result3996;
		result_out3997<=result3997;
		result_out3998<=result3998;
		result_out3999<=result3999;
		result_out4000<=result4000;
		result_out4001<=result4001;
		result_out4002<=result4002;
		result_out4003<=result4003;
		result_out4004<=result4004;
		result_out4005<=result4005;
		result_out4006<=result4006;
		result_out4007<=result4007;
		result_out4008<=result4008;
		result_out4009<=result4009;
		result_out4010<=result4010;
		result_out4011<=result4011;
		result_out4012<=result4012;
		result_out4013<=result4013;
		result_out4014<=result4014;
		result_out4015<=result4015;
		result_out4016<=result4016;
		result_out4017<=result4017;
		result_out4018<=result4018;
		result_out4019<=result4019;
		result_out4020<=result4020;
		result_out4021<=result4021;
		result_out4022<=result4022;
		result_out4023<=result4023;
		result_out4024<=result4024;
		result_out4025<=result4025;
		result_out4026<=result4026;
		result_out4027<=result4027;
		result_out4028<=result4028;
		result_out4029<=result4029;
		result_out4030<=result4030;
		result_out4031<=result4031;
		result_out4032<=result4032;
		result_out4033<=result4033;
		result_out4034<=result4034;
		result_out4035<=result4035;
		result_out4036<=result4036;
		result_out4037<=result4037;
		result_out4038<=result4038;
		result_out4039<=result4039;
		result_out4040<=result4040;
		result_out4041<=result4041;
		result_out4042<=result4042;
		result_out4043<=result4043;
		result_out4044<=result4044;
		result_out4045<=result4045;
		result_out4046<=result4046;
		result_out4047<=result4047;
		result_out4048<=result4048;
		result_out4049<=result4049;
		result_out4050<=result4050;
		result_out4051<=result4051;
		result_out4052<=result4052;
		result_out4053<=result4053;
		result_out4054<=result4054;
		result_out4055<=result4055;
		result_out4056<=result4056;
		result_out4057<=result4057;
		result_out4058<=result4058;
		result_out4059<=result4059;
		result_out4060<=result4060;
		result_out4061<=result4061;
		result_out4062<=result4062;
		result_out4063<=result4063;
		result_out4064<=result4064;
		result_out4065<=result4065;
		result_out4066<=result4066;
		result_out4067<=result4067;
		result_out4068<=result4068;
		result_out4069<=result4069;
		result_out4070<=result4070;
		result_out4071<=result4071;
		result_out4072<=result4072;
		result_out4073<=result4073;
		result_out4074<=result4074;
		result_out4075<=result4075;
		result_out4076<=result4076;
		result_out4077<=result4077;
		result_out4078<=result4078;
		result_out4079<=result4079;
		result_out4080<=result4080;
		result_out4081<=result4081;
		result_out4082<=result4082;
		result_out4083<=result4083;
		result_out4084<=result4084;
		result_out4085<=result4085;
		result_out4086<=result4086;
		result_out4087<=result4087;
		result_out4088<=result4088;
		result_out4089<=result4089;
		result_out4090<=result4090;
		result_out4091<=result4091;
		result_out4092<=result4092;
		result_out4093<=result4093;
		result_out4094<=result4094;
		result_out4095<=result4095;
		if(count == 190) begin
            done <= 1;
            count <= 0;
        end
        else begin
            done <= 0;
            count <= count + 1;
        end
    end
end
endmodule
