`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/19/2023 07:05:12 PM
// Design Name: 
// Module Name: sys_arr32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module syst_arr32(
	input [15:0] inp_w0,inp_w32,inp_w64,inp_w96,inp_w128,inp_w160,inp_w192,inp_w224,inp_w256,inp_w288,inp_w320,inp_w352,inp_w384,inp_w416,inp_w448,inp_w480,inp_w512,inp_w544,inp_w576,inp_w608,inp_w640,inp_w672,inp_w704,inp_w736,inp_w768,inp_w800,inp_w832,inp_w864,inp_w896,inp_w928,inp_w960,inp_w992,inp_n0,inp_n1,inp_n2,inp_n3,inp_n4,inp_n5,inp_n6,inp_n7,inp_n8,inp_n9,inp_n10,inp_n11,inp_n12,inp_n13,inp_n14,inp_n15,inp_n16,inp_n17,inp_n18,inp_n19,inp_n20,inp_n21,inp_n22,inp_n23,inp_n24,inp_n25,inp_n26,inp_n27,inp_n28,inp_n29,inp_n30,inp_n31,
	output reg [15:0]  result_out0, result_out1, result_out2, result_out3, result_out4, result_out5, result_out6, result_out7, result_out8, result_out9, result_out10, result_out11, result_out12, result_out13, result_out14, result_out15, result_out16, result_out17, result_out18, result_out19, result_out20, result_out21, result_out22, result_out23, result_out24, result_out25, result_out26, result_out27, result_out28, result_out29, result_out30, result_out31,result_out32, result_out33, result_out34, result_out35, result_out36, result_out37, result_out38, result_out39, result_out40, result_out41, result_out42, result_out43, result_out44, result_out45, result_out46, result_out47, result_out48, result_out49, result_out50, result_out51, result_out52, result_out53, result_out54, result_out55, result_out56, result_out57, result_out58, result_out59, result_out60, result_out61, result_out62, result_out63, result_out64, result_out65, result_out66, result_out67, result_out68, result_out69, result_out70, result_out71, result_out72, result_out73, result_out74, result_out75, result_out76, result_out77, result_out78, result_out79, result_out80, result_out81, result_out82, result_out83, result_out84, result_out85, result_out86, result_out87, result_out88, result_out89, result_out90, result_out91, result_out92, result_out93, result_out94, result_out95, result_out96, result_out97, result_out98, result_out99, result_out100, result_out101, result_out102, result_out103, result_out104, result_out105, result_out106, result_out107, result_out108, result_out109, result_out110, result_out111, result_out112, result_out113, result_out114, result_out115, result_out116, result_out117, result_out118, result_out119, result_out120, result_out121, result_out122, result_out123, result_out124, result_out125, result_out126, result_out127, result_out128, result_out129, result_out130, result_out131, result_out132, result_out133, result_out134, result_out135, result_out136, result_out137, result_out138, result_out139, result_out140, result_out141, result_out142, result_out143, result_out144, result_out145, result_out146, result_out147, result_out148, result_out149, result_out150, result_out151, result_out152, result_out153, result_out154, result_out155, result_out156, result_out157, result_out158, result_out159, result_out160, result_out161, result_out162, result_out163, result_out164, result_out165, result_out166, result_out167, result_out168, result_out169, result_out170, result_out171, result_out172, result_out173, result_out174, result_out175, result_out176, result_out177, result_out178, result_out179, result_out180, result_out181, result_out182, result_out183, result_out184, result_out185, result_out186, result_out187, result_out188, result_out189, result_out190, result_out191, result_out192, result_out193, result_out194, result_out195, result_out196, result_out197, result_out198, result_out199, result_out200, result_out201, result_out202, result_out203, result_out204, result_out205, result_out206, result_out207, result_out208, result_out209, result_out210, result_out211, result_out212, result_out213, result_out214, result_out215, result_out216, result_out217, result_out218, result_out219, result_out220, result_out221, result_out222, result_out223, result_out224, result_out225, result_out226, result_out227, result_out228, result_out229, result_out230, result_out231, result_out232, result_out233, result_out234, result_out235, result_out236, result_out237, result_out238, result_out239, result_out240, result_out241, result_out242, result_out243, result_out244, result_out245, result_out246, result_out247, result_out248, result_out249, result_out250, result_out251, result_out252, result_out253, result_out254, result_out255, result_out256, result_out257, result_out258, result_out259, result_out260, result_out261, result_out262, result_out263, result_out264, result_out265, result_out266, result_out267, result_out268, result_out269, result_out270, result_out271, result_out272, result_out273, result_out274, result_out275, result_out276, result_out277, result_out278, result_out279, result_out280, result_out281, result_out282, result_out283, result_out284, result_out285, result_out286, result_out287, result_out288, result_out289, result_out290, result_out291, result_out292, result_out293, result_out294, result_out295, result_out296, result_out297, result_out298, result_out299, result_out300, result_out301, result_out302, result_out303, result_out304, result_out305, result_out306, result_out307, result_out308, result_out309, result_out310, result_out311, result_out312, result_out313, result_out314, result_out315, result_out316, result_out317, result_out318, result_out319, result_out320, result_out321, result_out322, result_out323, result_out324, result_out325, result_out326, result_out327, result_out328, result_out329, result_out330, result_out331, result_out332, result_out333, result_out334, result_out335, result_out336, result_out337, result_out338, result_out339, result_out340, result_out341, result_out342, result_out343, result_out344, result_out345, result_out346, result_out347, result_out348, result_out349, result_out350, result_out351, result_out352, result_out353, result_out354, result_out355, result_out356, result_out357, result_out358, result_out359, result_out360, result_out361, result_out362, result_out363, result_out364, result_out365, result_out366, result_out367, result_out368, result_out369, result_out370, result_out371, result_out372, result_out373, result_out374, result_out375, result_out376, result_out377, result_out378, result_out379, result_out380, result_out381, result_out382, result_out383, result_out384, result_out385, result_out386, result_out387, result_out388, result_out389, result_out390, result_out391, result_out392, result_out393, result_out394, result_out395, result_out396, result_out397, result_out398, result_out399, result_out400, result_out401, result_out402, result_out403, result_out404, result_out405, result_out406, result_out407, result_out408, result_out409, result_out410, result_out411, result_out412, result_out413, result_out414, result_out415, result_out416, result_out417, result_out418, result_out419, result_out420, result_out421, result_out422, result_out423, result_out424, result_out425, result_out426, result_out427, result_out428, result_out429, result_out430, result_out431, result_out432, result_out433, result_out434, result_out435, result_out436, result_out437, result_out438, result_out439, result_out440, result_out441, result_out442, result_out443, result_out444, result_out445, result_out446, result_out447, result_out448, result_out449, result_out450, result_out451, result_out452, result_out453, result_out454, result_out455, result_out456, result_out457, result_out458, result_out459, result_out460, result_out461, result_out462, result_out463, result_out464, result_out465, result_out466, result_out467, result_out468, result_out469, result_out470, result_out471, result_out472, result_out473, result_out474, result_out475, result_out476, result_out477, result_out478, result_out479, result_out480, result_out481, result_out482, result_out483, result_out484, result_out485, result_out486, result_out487, result_out488, result_out489, result_out490, result_out491, result_out492, result_out493, result_out494, result_out495, result_out496, result_out497, result_out498, result_out499, result_out500, result_out501, result_out502, result_out503, result_out504, result_out505, result_out506, result_out507, result_out508, result_out509, result_out510, result_out511, result_out512, result_out513, result_out514, result_out515, result_out516, result_out517, result_out518, result_out519, result_out520, result_out521, result_out522, result_out523, result_out524, result_out525, result_out526, result_out527, result_out528, result_out529, result_out530, result_out531, result_out532, result_out533, result_out534, result_out535, result_out536, result_out537, result_out538, result_out539, result_out540, result_out541, result_out542, result_out543, result_out544, result_out545, result_out546, result_out547, result_out548, result_out549, result_out550, result_out551, result_out552, result_out553, result_out554, result_out555, result_out556, result_out557, result_out558, result_out559, result_out560, result_out561, result_out562, result_out563, result_out564, result_out565, result_out566, result_out567, result_out568, result_out569, result_out570, result_out571, result_out572, result_out573, result_out574, result_out575, result_out576, result_out577, result_out578, result_out579, result_out580, result_out581, result_out582, result_out583, result_out584, result_out585, result_out586, result_out587, result_out588, result_out589, result_out590, result_out591, result_out592, result_out593, result_out594, result_out595, result_out596, result_out597, result_out598, result_out599, result_out600, result_out601, result_out602, result_out603, result_out604, result_out605, result_out606, result_out607, result_out608, result_out609, result_out610, result_out611, result_out612, result_out613, result_out614, result_out615, result_out616, result_out617, result_out618, result_out619, result_out620, result_out621, result_out622, result_out623, result_out624, result_out625, result_out626, result_out627, result_out628, result_out629, result_out630, result_out631, result_out632, result_out633, result_out634, result_out635, result_out636, result_out637, result_out638, result_out639, result_out640, result_out641, result_out642, result_out643, result_out644, result_out645, result_out646, result_out647, result_out648, result_out649, result_out650, result_out651, result_out652, result_out653, result_out654, result_out655, result_out656, result_out657, result_out658, result_out659, result_out660, result_out661, result_out662, result_out663, result_out664, result_out665, result_out666, result_out667, result_out668, result_out669, result_out670, result_out671, result_out672, result_out673, result_out674, result_out675, result_out676, result_out677, result_out678, result_out679, result_out680, result_out681, result_out682, result_out683, result_out684, result_out685, result_out686, result_out687, result_out688, result_out689, result_out690, result_out691, result_out692, result_out693, result_out694, result_out695, result_out696, result_out697, result_out698, result_out699, result_out700, result_out701, result_out702, result_out703, result_out704, result_out705, result_out706, result_out707, result_out708, result_out709, result_out710, result_out711, result_out712, result_out713, result_out714, result_out715, result_out716, result_out717, result_out718, result_out719, result_out720, result_out721, result_out722, result_out723, result_out724, result_out725, result_out726, result_out727, result_out728, result_out729, result_out730, result_out731, result_out732, result_out733, result_out734, result_out735, result_out736, result_out737, result_out738, result_out739, result_out740, result_out741, result_out742, result_out743, result_out744, result_out745, result_out746, result_out747, result_out748, result_out749, result_out750, result_out751, result_out752, result_out753, result_out754, result_out755, result_out756, result_out757, result_out758, result_out759, result_out760, result_out761, result_out762, result_out763, result_out764, result_out765, result_out766, result_out767, result_out768, result_out769, result_out770, result_out771, result_out772, result_out773, result_out774, result_out775, result_out776, result_out777, result_out778, result_out779, result_out780, result_out781, result_out782, result_out783, result_out784, result_out785, result_out786, result_out787, result_out788, result_out789, result_out790, result_out791, result_out792, result_out793, result_out794, result_out795, result_out796, result_out797, result_out798, result_out799, result_out800, result_out801, result_out802, result_out803, result_out804, result_out805, result_out806, result_out807, result_out808, result_out809, result_out810, result_out811, result_out812, result_out813, result_out814, result_out815, result_out816, result_out817, result_out818, result_out819, result_out820, result_out821, result_out822, result_out823, result_out824, result_out825, result_out826, result_out827, result_out828, result_out829, result_out830, result_out831, result_out832, result_out833, result_out834, result_out835, result_out836, result_out837, result_out838, result_out839, result_out840, result_out841, result_out842, result_out843, result_out844, result_out845, result_out846, result_out847, result_out848, result_out849, result_out850, result_out851, result_out852, result_out853, result_out854, result_out855, result_out856, result_out857, result_out858, result_out859, result_out860, result_out861, result_out862, result_out863, result_out864, result_out865, result_out866, result_out867, result_out868, result_out869, result_out870, result_out871, result_out872, result_out873, result_out874, result_out875, result_out876, result_out877, result_out878, result_out879, result_out880, result_out881, result_out882, result_out883, result_out884, result_out885, result_out886, result_out887, result_out888, result_out889, result_out890, result_out891, result_out892, result_out893, result_out894, result_out895, result_out896, result_out897, result_out898, result_out899, result_out900, result_out901, result_out902, result_out903, result_out904, result_out905, result_out906, result_out907, result_out908, result_out909, result_out910, result_out911, result_out912, result_out913, result_out914, result_out915, result_out916, result_out917, result_out918, result_out919, result_out920, result_out921, result_out922, result_out923, result_out924, result_out925, result_out926, result_out927, result_out928, result_out929, result_out930, result_out931, result_out932, result_out933, result_out934, result_out935, result_out936, result_out937, result_out938, result_out939, result_out940, result_out941, result_out942, result_out943, result_out944, result_out945, result_out946, result_out947, result_out948, result_out949, result_out950, result_out951, result_out952, result_out953, result_out954, result_out955, result_out956, result_out957, result_out958, result_out959, result_out960, result_out961, result_out962, result_out963, result_out964, result_out965, result_out966, result_out967, result_out968, result_out969, result_out970, result_out971, result_out972, result_out973, result_out974, result_out975, result_out976, result_out977, result_out978, result_out979, result_out980, result_out981, result_out982, result_out983, result_out984, result_out985, result_out986, result_out987, result_out988, result_out989, result_out990, result_out991, result_out992, result_out993, result_out994, result_out995, result_out996, result_out997, result_out998, result_out999, result_out1000, result_out1001, result_out1002, result_out1003, result_out1004, result_out1005, result_out1006, result_out1007, result_out1008, result_out1009, result_out1010, result_out1011, result_out1012, result_out1013, result_out1014, result_out1015, result_out1016, result_out1017, result_out1018, result_out1019, result_out1020, result_out1021, result_out1022, result_out1023, 
	output reg done,
	input clk,rst
); 

reg [6:0] count;

wire  [15:0] out_s0;
wire  [15:0] out_s1;
wire  [15:0] out_s2;
wire  [15:0] out_s3;
wire  [15:0] out_s4;
wire  [15:0] out_s5;
wire  [15:0] out_s6;
wire  [15:0] out_s7;
wire  [15:0] out_s8;
wire  [15:0] out_s9;
wire  [15:0] out_s10;
wire  [15:0] out_s11;
wire  [15:0] out_s12;
wire  [15:0] out_s13;
wire  [15:0] out_s14;
wire  [15:0] out_s15;
wire  [15:0] out_s16;
wire  [15:0] out_s17;
wire  [15:0] out_s18;
wire  [15:0] out_s19;
wire  [15:0] out_s20;
wire  [15:0] out_s21;
wire  [15:0] out_s22;
wire  [15:0] out_s23;
wire  [15:0] out_s24;
wire  [15:0] out_s25;
wire  [15:0] out_s26;
wire  [15:0] out_s27;
wire  [15:0] out_s28;
wire  [15:0] out_s29;
wire  [15:0] out_s30;
wire  [15:0] out_s31;
wire  [15:0] out_s32;
wire  [15:0] out_s33;
wire  [15:0] out_s34;
wire  [15:0] out_s35;
wire  [15:0] out_s36;
wire  [15:0] out_s37;
wire  [15:0] out_s38;
wire  [15:0] out_s39;
wire  [15:0] out_s40;
wire  [15:0] out_s41;
wire  [15:0] out_s42;
wire  [15:0] out_s43;
wire  [15:0] out_s44;
wire  [15:0] out_s45;
wire  [15:0] out_s46;
wire  [15:0] out_s47;
wire  [15:0] out_s48;
wire  [15:0] out_s49;
wire  [15:0] out_s50;
wire  [15:0] out_s51;
wire  [15:0] out_s52;
wire  [15:0] out_s53;
wire  [15:0] out_s54;
wire  [15:0] out_s55;
wire  [15:0] out_s56;
wire  [15:0] out_s57;
wire  [15:0] out_s58;
wire  [15:0] out_s59;
wire  [15:0] out_s60;
wire  [15:0] out_s61;
wire  [15:0] out_s62;
wire  [15:0] out_s63;
wire  [15:0] out_s64;
wire  [15:0] out_s65;
wire  [15:0] out_s66;
wire  [15:0] out_s67;
wire  [15:0] out_s68;
wire  [15:0] out_s69;
wire  [15:0] out_s70;
wire  [15:0] out_s71;
wire  [15:0] out_s72;
wire  [15:0] out_s73;
wire  [15:0] out_s74;
wire  [15:0] out_s75;
wire  [15:0] out_s76;
wire  [15:0] out_s77;
wire  [15:0] out_s78;
wire  [15:0] out_s79;
wire  [15:0] out_s80;
wire  [15:0] out_s81;
wire  [15:0] out_s82;
wire  [15:0] out_s83;
wire  [15:0] out_s84;
wire  [15:0] out_s85;
wire  [15:0] out_s86;
wire  [15:0] out_s87;
wire  [15:0] out_s88;
wire  [15:0] out_s89;
wire  [15:0] out_s90;
wire  [15:0] out_s91;
wire  [15:0] out_s92;
wire  [15:0] out_s93;
wire  [15:0] out_s94;
wire  [15:0] out_s95;
wire  [15:0] out_s96;
wire  [15:0] out_s97;
wire  [15:0] out_s98;
wire  [15:0] out_s99;
wire  [15:0] out_s100;
wire  [15:0] out_s101;
wire  [15:0] out_s102;
wire  [15:0] out_s103;
wire  [15:0] out_s104;
wire  [15:0] out_s105;
wire  [15:0] out_s106;
wire  [15:0] out_s107;
wire  [15:0] out_s108;
wire  [15:0] out_s109;
wire  [15:0] out_s110;
wire  [15:0] out_s111;
wire  [15:0] out_s112;
wire  [15:0] out_s113;
wire  [15:0] out_s114;
wire  [15:0] out_s115;
wire  [15:0] out_s116;
wire  [15:0] out_s117;
wire  [15:0] out_s118;
wire  [15:0] out_s119;
wire  [15:0] out_s120;
wire  [15:0] out_s121;
wire  [15:0] out_s122;
wire  [15:0] out_s123;
wire  [15:0] out_s124;
wire  [15:0] out_s125;
wire  [15:0] out_s126;
wire  [15:0] out_s127;
wire  [15:0] out_s128;
wire  [15:0] out_s129;
wire  [15:0] out_s130;
wire  [15:0] out_s131;
wire  [15:0] out_s132;
wire  [15:0] out_s133;
wire  [15:0] out_s134;
wire  [15:0] out_s135;
wire  [15:0] out_s136;
wire  [15:0] out_s137;
wire  [15:0] out_s138;
wire  [15:0] out_s139;
wire  [15:0] out_s140;
wire  [15:0] out_s141;
wire  [15:0] out_s142;
wire  [15:0] out_s143;
wire  [15:0] out_s144;
wire  [15:0] out_s145;
wire  [15:0] out_s146;
wire  [15:0] out_s147;
wire  [15:0] out_s148;
wire  [15:0] out_s149;
wire  [15:0] out_s150;
wire  [15:0] out_s151;
wire  [15:0] out_s152;
wire  [15:0] out_s153;
wire  [15:0] out_s154;
wire  [15:0] out_s155;
wire  [15:0] out_s156;
wire  [15:0] out_s157;
wire  [15:0] out_s158;
wire  [15:0] out_s159;
wire  [15:0] out_s160;
wire  [15:0] out_s161;
wire  [15:0] out_s162;
wire  [15:0] out_s163;
wire  [15:0] out_s164;
wire  [15:0] out_s165;
wire  [15:0] out_s166;
wire  [15:0] out_s167;
wire  [15:0] out_s168;
wire  [15:0] out_s169;
wire  [15:0] out_s170;
wire  [15:0] out_s171;
wire  [15:0] out_s172;
wire  [15:0] out_s173;
wire  [15:0] out_s174;
wire  [15:0] out_s175;
wire  [15:0] out_s176;
wire  [15:0] out_s177;
wire  [15:0] out_s178;
wire  [15:0] out_s179;
wire  [15:0] out_s180;
wire  [15:0] out_s181;
wire  [15:0] out_s182;
wire  [15:0] out_s183;
wire  [15:0] out_s184;
wire  [15:0] out_s185;
wire  [15:0] out_s186;
wire  [15:0] out_s187;
wire  [15:0] out_s188;
wire  [15:0] out_s189;
wire  [15:0] out_s190;
wire  [15:0] out_s191;
wire  [15:0] out_s192;
wire  [15:0] out_s193;
wire  [15:0] out_s194;
wire  [15:0] out_s195;
wire  [15:0] out_s196;
wire  [15:0] out_s197;
wire  [15:0] out_s198;
wire  [15:0] out_s199;
wire  [15:0] out_s200;
wire  [15:0] out_s201;
wire  [15:0] out_s202;
wire  [15:0] out_s203;
wire  [15:0] out_s204;
wire  [15:0] out_s205;
wire  [15:0] out_s206;
wire  [15:0] out_s207;
wire  [15:0] out_s208;
wire  [15:0] out_s209;
wire  [15:0] out_s210;
wire  [15:0] out_s211;
wire  [15:0] out_s212;
wire  [15:0] out_s213;
wire  [15:0] out_s214;
wire  [15:0] out_s215;
wire  [15:0] out_s216;
wire  [15:0] out_s217;
wire  [15:0] out_s218;
wire  [15:0] out_s219;
wire  [15:0] out_s220;
wire  [15:0] out_s221;
wire  [15:0] out_s222;
wire  [15:0] out_s223;
wire  [15:0] out_s224;
wire  [15:0] out_s225;
wire  [15:0] out_s226;
wire  [15:0] out_s227;
wire  [15:0] out_s228;
wire  [15:0] out_s229;
wire  [15:0] out_s230;
wire  [15:0] out_s231;
wire  [15:0] out_s232;
wire  [15:0] out_s233;
wire  [15:0] out_s234;
wire  [15:0] out_s235;
wire  [15:0] out_s236;
wire  [15:0] out_s237;
wire  [15:0] out_s238;
wire  [15:0] out_s239;
wire  [15:0] out_s240;
wire  [15:0] out_s241;
wire  [15:0] out_s242;
wire  [15:0] out_s243;
wire  [15:0] out_s244;
wire  [15:0] out_s245;
wire  [15:0] out_s246;
wire  [15:0] out_s247;
wire  [15:0] out_s248;
wire  [15:0] out_s249;
wire  [15:0] out_s250;
wire  [15:0] out_s251;
wire  [15:0] out_s252;
wire  [15:0] out_s253;
wire  [15:0] out_s254;
wire  [15:0] out_s255;
wire  [15:0] out_s256;
wire  [15:0] out_s257;
wire  [15:0] out_s258;
wire  [15:0] out_s259;
wire  [15:0] out_s260;
wire  [15:0] out_s261;
wire  [15:0] out_s262;
wire  [15:0] out_s263;
wire  [15:0] out_s264;
wire  [15:0] out_s265;
wire  [15:0] out_s266;
wire  [15:0] out_s267;
wire  [15:0] out_s268;
wire  [15:0] out_s269;
wire  [15:0] out_s270;
wire  [15:0] out_s271;
wire  [15:0] out_s272;
wire  [15:0] out_s273;
wire  [15:0] out_s274;
wire  [15:0] out_s275;
wire  [15:0] out_s276;
wire  [15:0] out_s277;
wire  [15:0] out_s278;
wire  [15:0] out_s279;
wire  [15:0] out_s280;
wire  [15:0] out_s281;
wire  [15:0] out_s282;
wire  [15:0] out_s283;
wire  [15:0] out_s284;
wire  [15:0] out_s285;
wire  [15:0] out_s286;
wire  [15:0] out_s287;
wire  [15:0] out_s288;
wire  [15:0] out_s289;
wire  [15:0] out_s290;
wire  [15:0] out_s291;
wire  [15:0] out_s292;
wire  [15:0] out_s293;
wire  [15:0] out_s294;
wire  [15:0] out_s295;
wire  [15:0] out_s296;
wire  [15:0] out_s297;
wire  [15:0] out_s298;
wire  [15:0] out_s299;
wire  [15:0] out_s300;
wire  [15:0] out_s301;
wire  [15:0] out_s302;
wire  [15:0] out_s303;
wire  [15:0] out_s304;
wire  [15:0] out_s305;
wire  [15:0] out_s306;
wire  [15:0] out_s307;
wire  [15:0] out_s308;
wire  [15:0] out_s309;
wire  [15:0] out_s310;
wire  [15:0] out_s311;
wire  [15:0] out_s312;
wire  [15:0] out_s313;
wire  [15:0] out_s314;
wire  [15:0] out_s315;
wire  [15:0] out_s316;
wire  [15:0] out_s317;
wire  [15:0] out_s318;
wire  [15:0] out_s319;
wire  [15:0] out_s320;
wire  [15:0] out_s321;
wire  [15:0] out_s322;
wire  [15:0] out_s323;
wire  [15:0] out_s324;
wire  [15:0] out_s325;
wire  [15:0] out_s326;
wire  [15:0] out_s327;
wire  [15:0] out_s328;
wire  [15:0] out_s329;
wire  [15:0] out_s330;
wire  [15:0] out_s331;
wire  [15:0] out_s332;
wire  [15:0] out_s333;
wire  [15:0] out_s334;
wire  [15:0] out_s335;
wire  [15:0] out_s336;
wire  [15:0] out_s337;
wire  [15:0] out_s338;
wire  [15:0] out_s339;
wire  [15:0] out_s340;
wire  [15:0] out_s341;
wire  [15:0] out_s342;
wire  [15:0] out_s343;
wire  [15:0] out_s344;
wire  [15:0] out_s345;
wire  [15:0] out_s346;
wire  [15:0] out_s347;
wire  [15:0] out_s348;
wire  [15:0] out_s349;
wire  [15:0] out_s350;
wire  [15:0] out_s351;
wire  [15:0] out_s352;
wire  [15:0] out_s353;
wire  [15:0] out_s354;
wire  [15:0] out_s355;
wire  [15:0] out_s356;
wire  [15:0] out_s357;
wire  [15:0] out_s358;
wire  [15:0] out_s359;
wire  [15:0] out_s360;
wire  [15:0] out_s361;
wire  [15:0] out_s362;
wire  [15:0] out_s363;
wire  [15:0] out_s364;
wire  [15:0] out_s365;
wire  [15:0] out_s366;
wire  [15:0] out_s367;
wire  [15:0] out_s368;
wire  [15:0] out_s369;
wire  [15:0] out_s370;
wire  [15:0] out_s371;
wire  [15:0] out_s372;
wire  [15:0] out_s373;
wire  [15:0] out_s374;
wire  [15:0] out_s375;
wire  [15:0] out_s376;
wire  [15:0] out_s377;
wire  [15:0] out_s378;
wire  [15:0] out_s379;
wire  [15:0] out_s380;
wire  [15:0] out_s381;
wire  [15:0] out_s382;
wire  [15:0] out_s383;
wire  [15:0] out_s384;
wire  [15:0] out_s385;
wire  [15:0] out_s386;
wire  [15:0] out_s387;
wire  [15:0] out_s388;
wire  [15:0] out_s389;
wire  [15:0] out_s390;
wire  [15:0] out_s391;
wire  [15:0] out_s392;
wire  [15:0] out_s393;
wire  [15:0] out_s394;
wire  [15:0] out_s395;
wire  [15:0] out_s396;
wire  [15:0] out_s397;
wire  [15:0] out_s398;
wire  [15:0] out_s399;
wire  [15:0] out_s400;
wire  [15:0] out_s401;
wire  [15:0] out_s402;
wire  [15:0] out_s403;
wire  [15:0] out_s404;
wire  [15:0] out_s405;
wire  [15:0] out_s406;
wire  [15:0] out_s407;
wire  [15:0] out_s408;
wire  [15:0] out_s409;
wire  [15:0] out_s410;
wire  [15:0] out_s411;
wire  [15:0] out_s412;
wire  [15:0] out_s413;
wire  [15:0] out_s414;
wire  [15:0] out_s415;
wire  [15:0] out_s416;
wire  [15:0] out_s417;
wire  [15:0] out_s418;
wire  [15:0] out_s419;
wire  [15:0] out_s420;
wire  [15:0] out_s421;
wire  [15:0] out_s422;
wire  [15:0] out_s423;
wire  [15:0] out_s424;
wire  [15:0] out_s425;
wire  [15:0] out_s426;
wire  [15:0] out_s427;
wire  [15:0] out_s428;
wire  [15:0] out_s429;
wire  [15:0] out_s430;
wire  [15:0] out_s431;
wire  [15:0] out_s432;
wire  [15:0] out_s433;
wire  [15:0] out_s434;
wire  [15:0] out_s435;
wire  [15:0] out_s436;
wire  [15:0] out_s437;
wire  [15:0] out_s438;
wire  [15:0] out_s439;
wire  [15:0] out_s440;
wire  [15:0] out_s441;
wire  [15:0] out_s442;
wire  [15:0] out_s443;
wire  [15:0] out_s444;
wire  [15:0] out_s445;
wire  [15:0] out_s446;
wire  [15:0] out_s447;
wire  [15:0] out_s448;
wire  [15:0] out_s449;
wire  [15:0] out_s450;
wire  [15:0] out_s451;
wire  [15:0] out_s452;
wire  [15:0] out_s453;
wire  [15:0] out_s454;
wire  [15:0] out_s455;
wire  [15:0] out_s456;
wire  [15:0] out_s457;
wire  [15:0] out_s458;
wire  [15:0] out_s459;
wire  [15:0] out_s460;
wire  [15:0] out_s461;
wire  [15:0] out_s462;
wire  [15:0] out_s463;
wire  [15:0] out_s464;
wire  [15:0] out_s465;
wire  [15:0] out_s466;
wire  [15:0] out_s467;
wire  [15:0] out_s468;
wire  [15:0] out_s469;
wire  [15:0] out_s470;
wire  [15:0] out_s471;
wire  [15:0] out_s472;
wire  [15:0] out_s473;
wire  [15:0] out_s474;
wire  [15:0] out_s475;
wire  [15:0] out_s476;
wire  [15:0] out_s477;
wire  [15:0] out_s478;
wire  [15:0] out_s479;
wire  [15:0] out_s480;
wire  [15:0] out_s481;
wire  [15:0] out_s482;
wire  [15:0] out_s483;
wire  [15:0] out_s484;
wire  [15:0] out_s485;
wire  [15:0] out_s486;
wire  [15:0] out_s487;
wire  [15:0] out_s488;
wire  [15:0] out_s489;
wire  [15:0] out_s490;
wire  [15:0] out_s491;
wire  [15:0] out_s492;
wire  [15:0] out_s493;
wire  [15:0] out_s494;
wire  [15:0] out_s495;
wire  [15:0] out_s496;
wire  [15:0] out_s497;
wire  [15:0] out_s498;
wire  [15:0] out_s499;
wire  [15:0] out_s500;
wire  [15:0] out_s501;
wire  [15:0] out_s502;
wire  [15:0] out_s503;
wire  [15:0] out_s504;
wire  [15:0] out_s505;
wire  [15:0] out_s506;
wire  [15:0] out_s507;
wire  [15:0] out_s508;
wire  [15:0] out_s509;
wire  [15:0] out_s510;
wire  [15:0] out_s511;
wire  [15:0] out_s512;
wire  [15:0] out_s513;
wire  [15:0] out_s514;
wire  [15:0] out_s515;
wire  [15:0] out_s516;
wire  [15:0] out_s517;
wire  [15:0] out_s518;
wire  [15:0] out_s519;
wire  [15:0] out_s520;
wire  [15:0] out_s521;
wire  [15:0] out_s522;
wire  [15:0] out_s523;
wire  [15:0] out_s524;
wire  [15:0] out_s525;
wire  [15:0] out_s526;
wire  [15:0] out_s527;
wire  [15:0] out_s528;
wire  [15:0] out_s529;
wire  [15:0] out_s530;
wire  [15:0] out_s531;
wire  [15:0] out_s532;
wire  [15:0] out_s533;
wire  [15:0] out_s534;
wire  [15:0] out_s535;
wire  [15:0] out_s536;
wire  [15:0] out_s537;
wire  [15:0] out_s538;
wire  [15:0] out_s539;
wire  [15:0] out_s540;
wire  [15:0] out_s541;
wire  [15:0] out_s542;
wire  [15:0] out_s543;
wire  [15:0] out_s544;
wire  [15:0] out_s545;
wire  [15:0] out_s546;
wire  [15:0] out_s547;
wire  [15:0] out_s548;
wire  [15:0] out_s549;
wire  [15:0] out_s550;
wire  [15:0] out_s551;
wire  [15:0] out_s552;
wire  [15:0] out_s553;
wire  [15:0] out_s554;
wire  [15:0] out_s555;
wire  [15:0] out_s556;
wire  [15:0] out_s557;
wire  [15:0] out_s558;
wire  [15:0] out_s559;
wire  [15:0] out_s560;
wire  [15:0] out_s561;
wire  [15:0] out_s562;
wire  [15:0] out_s563;
wire  [15:0] out_s564;
wire  [15:0] out_s565;
wire  [15:0] out_s566;
wire  [15:0] out_s567;
wire  [15:0] out_s568;
wire  [15:0] out_s569;
wire  [15:0] out_s570;
wire  [15:0] out_s571;
wire  [15:0] out_s572;
wire  [15:0] out_s573;
wire  [15:0] out_s574;
wire  [15:0] out_s575;
wire  [15:0] out_s576;
wire  [15:0] out_s577;
wire  [15:0] out_s578;
wire  [15:0] out_s579;
wire  [15:0] out_s580;
wire  [15:0] out_s581;
wire  [15:0] out_s582;
wire  [15:0] out_s583;
wire  [15:0] out_s584;
wire  [15:0] out_s585;
wire  [15:0] out_s586;
wire  [15:0] out_s587;
wire  [15:0] out_s588;
wire  [15:0] out_s589;
wire  [15:0] out_s590;
wire  [15:0] out_s591;
wire  [15:0] out_s592;
wire  [15:0] out_s593;
wire  [15:0] out_s594;
wire  [15:0] out_s595;
wire  [15:0] out_s596;
wire  [15:0] out_s597;
wire  [15:0] out_s598;
wire  [15:0] out_s599;
wire  [15:0] out_s600;
wire  [15:0] out_s601;
wire  [15:0] out_s602;
wire  [15:0] out_s603;
wire  [15:0] out_s604;
wire  [15:0] out_s605;
wire  [15:0] out_s606;
wire  [15:0] out_s607;
wire  [15:0] out_s608;
wire  [15:0] out_s609;
wire  [15:0] out_s610;
wire  [15:0] out_s611;
wire  [15:0] out_s612;
wire  [15:0] out_s613;
wire  [15:0] out_s614;
wire  [15:0] out_s615;
wire  [15:0] out_s616;
wire  [15:0] out_s617;
wire  [15:0] out_s618;
wire  [15:0] out_s619;
wire  [15:0] out_s620;
wire  [15:0] out_s621;
wire  [15:0] out_s622;
wire  [15:0] out_s623;
wire  [15:0] out_s624;
wire  [15:0] out_s625;
wire  [15:0] out_s626;
wire  [15:0] out_s627;
wire  [15:0] out_s628;
wire  [15:0] out_s629;
wire  [15:0] out_s630;
wire  [15:0] out_s631;
wire  [15:0] out_s632;
wire  [15:0] out_s633;
wire  [15:0] out_s634;
wire  [15:0] out_s635;
wire  [15:0] out_s636;
wire  [15:0] out_s637;
wire  [15:0] out_s638;
wire  [15:0] out_s639;
wire  [15:0] out_s640;
wire  [15:0] out_s641;
wire  [15:0] out_s642;
wire  [15:0] out_s643;
wire  [15:0] out_s644;
wire  [15:0] out_s645;
wire  [15:0] out_s646;
wire  [15:0] out_s647;
wire  [15:0] out_s648;
wire  [15:0] out_s649;
wire  [15:0] out_s650;
wire  [15:0] out_s651;
wire  [15:0] out_s652;
wire  [15:0] out_s653;
wire  [15:0] out_s654;
wire  [15:0] out_s655;
wire  [15:0] out_s656;
wire  [15:0] out_s657;
wire  [15:0] out_s658;
wire  [15:0] out_s659;
wire  [15:0] out_s660;
wire  [15:0] out_s661;
wire  [15:0] out_s662;
wire  [15:0] out_s663;
wire  [15:0] out_s664;
wire  [15:0] out_s665;
wire  [15:0] out_s666;
wire  [15:0] out_s667;
wire  [15:0] out_s668;
wire  [15:0] out_s669;
wire  [15:0] out_s670;
wire  [15:0] out_s671;
wire  [15:0] out_s672;
wire  [15:0] out_s673;
wire  [15:0] out_s674;
wire  [15:0] out_s675;
wire  [15:0] out_s676;
wire  [15:0] out_s677;
wire  [15:0] out_s678;
wire  [15:0] out_s679;
wire  [15:0] out_s680;
wire  [15:0] out_s681;
wire  [15:0] out_s682;
wire  [15:0] out_s683;
wire  [15:0] out_s684;
wire  [15:0] out_s685;
wire  [15:0] out_s686;
wire  [15:0] out_s687;
wire  [15:0] out_s688;
wire  [15:0] out_s689;
wire  [15:0] out_s690;
wire  [15:0] out_s691;
wire  [15:0] out_s692;
wire  [15:0] out_s693;
wire  [15:0] out_s694;
wire  [15:0] out_s695;
wire  [15:0] out_s696;
wire  [15:0] out_s697;
wire  [15:0] out_s698;
wire  [15:0] out_s699;
wire  [15:0] out_s700;
wire  [15:0] out_s701;
wire  [15:0] out_s702;
wire  [15:0] out_s703;
wire  [15:0] out_s704;
wire  [15:0] out_s705;
wire  [15:0] out_s706;
wire  [15:0] out_s707;
wire  [15:0] out_s708;
wire  [15:0] out_s709;
wire  [15:0] out_s710;
wire  [15:0] out_s711;
wire  [15:0] out_s712;
wire  [15:0] out_s713;
wire  [15:0] out_s714;
wire  [15:0] out_s715;
wire  [15:0] out_s716;
wire  [15:0] out_s717;
wire  [15:0] out_s718;
wire  [15:0] out_s719;
wire  [15:0] out_s720;
wire  [15:0] out_s721;
wire  [15:0] out_s722;
wire  [15:0] out_s723;
wire  [15:0] out_s724;
wire  [15:0] out_s725;
wire  [15:0] out_s726;
wire  [15:0] out_s727;
wire  [15:0] out_s728;
wire  [15:0] out_s729;
wire  [15:0] out_s730;
wire  [15:0] out_s731;
wire  [15:0] out_s732;
wire  [15:0] out_s733;
wire  [15:0] out_s734;
wire  [15:0] out_s735;
wire  [15:0] out_s736;
wire  [15:0] out_s737;
wire  [15:0] out_s738;
wire  [15:0] out_s739;
wire  [15:0] out_s740;
wire  [15:0] out_s741;
wire  [15:0] out_s742;
wire  [15:0] out_s743;
wire  [15:0] out_s744;
wire  [15:0] out_s745;
wire  [15:0] out_s746;
wire  [15:0] out_s747;
wire  [15:0] out_s748;
wire  [15:0] out_s749;
wire  [15:0] out_s750;
wire  [15:0] out_s751;
wire  [15:0] out_s752;
wire  [15:0] out_s753;
wire  [15:0] out_s754;
wire  [15:0] out_s755;
wire  [15:0] out_s756;
wire  [15:0] out_s757;
wire  [15:0] out_s758;
wire  [15:0] out_s759;
wire  [15:0] out_s760;
wire  [15:0] out_s761;
wire  [15:0] out_s762;
wire  [15:0] out_s763;
wire  [15:0] out_s764;
wire  [15:0] out_s765;
wire  [15:0] out_s766;
wire  [15:0] out_s767;
wire  [15:0] out_s768;
wire  [15:0] out_s769;
wire  [15:0] out_s770;
wire  [15:0] out_s771;
wire  [15:0] out_s772;
wire  [15:0] out_s773;
wire  [15:0] out_s774;
wire  [15:0] out_s775;
wire  [15:0] out_s776;
wire  [15:0] out_s777;
wire  [15:0] out_s778;
wire  [15:0] out_s779;
wire  [15:0] out_s780;
wire  [15:0] out_s781;
wire  [15:0] out_s782;
wire  [15:0] out_s783;
wire  [15:0] out_s784;
wire  [15:0] out_s785;
wire  [15:0] out_s786;
wire  [15:0] out_s787;
wire  [15:0] out_s788;
wire  [15:0] out_s789;
wire  [15:0] out_s790;
wire  [15:0] out_s791;
wire  [15:0] out_s792;
wire  [15:0] out_s793;
wire  [15:0] out_s794;
wire  [15:0] out_s795;
wire  [15:0] out_s796;
wire  [15:0] out_s797;
wire  [15:0] out_s798;
wire  [15:0] out_s799;
wire  [15:0] out_s800;
wire  [15:0] out_s801;
wire  [15:0] out_s802;
wire  [15:0] out_s803;
wire  [15:0] out_s804;
wire  [15:0] out_s805;
wire  [15:0] out_s806;
wire  [15:0] out_s807;
wire  [15:0] out_s808;
wire  [15:0] out_s809;
wire  [15:0] out_s810;
wire  [15:0] out_s811;
wire  [15:0] out_s812;
wire  [15:0] out_s813;
wire  [15:0] out_s814;
wire  [15:0] out_s815;
wire  [15:0] out_s816;
wire  [15:0] out_s817;
wire  [15:0] out_s818;
wire  [15:0] out_s819;
wire  [15:0] out_s820;
wire  [15:0] out_s821;
wire  [15:0] out_s822;
wire  [15:0] out_s823;
wire  [15:0] out_s824;
wire  [15:0] out_s825;
wire  [15:0] out_s826;
wire  [15:0] out_s827;
wire  [15:0] out_s828;
wire  [15:0] out_s829;
wire  [15:0] out_s830;
wire  [15:0] out_s831;
wire  [15:0] out_s832;
wire  [15:0] out_s833;
wire  [15:0] out_s834;
wire  [15:0] out_s835;
wire  [15:0] out_s836;
wire  [15:0] out_s837;
wire  [15:0] out_s838;
wire  [15:0] out_s839;
wire  [15:0] out_s840;
wire  [15:0] out_s841;
wire  [15:0] out_s842;
wire  [15:0] out_s843;
wire  [15:0] out_s844;
wire  [15:0] out_s845;
wire  [15:0] out_s846;
wire  [15:0] out_s847;
wire  [15:0] out_s848;
wire  [15:0] out_s849;
wire  [15:0] out_s850;
wire  [15:0] out_s851;
wire  [15:0] out_s852;
wire  [15:0] out_s853;
wire  [15:0] out_s854;
wire  [15:0] out_s855;
wire  [15:0] out_s856;
wire  [15:0] out_s857;
wire  [15:0] out_s858;
wire  [15:0] out_s859;
wire  [15:0] out_s860;
wire  [15:0] out_s861;
wire  [15:0] out_s862;
wire  [15:0] out_s863;
wire  [15:0] out_s864;
wire  [15:0] out_s865;
wire  [15:0] out_s866;
wire  [15:0] out_s867;
wire  [15:0] out_s868;
wire  [15:0] out_s869;
wire  [15:0] out_s870;
wire  [15:0] out_s871;
wire  [15:0] out_s872;
wire  [15:0] out_s873;
wire  [15:0] out_s874;
wire  [15:0] out_s875;
wire  [15:0] out_s876;
wire  [15:0] out_s877;
wire  [15:0] out_s878;
wire  [15:0] out_s879;
wire  [15:0] out_s880;
wire  [15:0] out_s881;
wire  [15:0] out_s882;
wire  [15:0] out_s883;
wire  [15:0] out_s884;
wire  [15:0] out_s885;
wire  [15:0] out_s886;
wire  [15:0] out_s887;
wire  [15:0] out_s888;
wire  [15:0] out_s889;
wire  [15:0] out_s890;
wire  [15:0] out_s891;
wire  [15:0] out_s892;
wire  [15:0] out_s893;
wire  [15:0] out_s894;
wire  [15:0] out_s895;
wire  [15:0] out_s896;
wire  [15:0] out_s897;
wire  [15:0] out_s898;
wire  [15:0] out_s899;
wire  [15:0] out_s900;
wire  [15:0] out_s901;
wire  [15:0] out_s902;
wire  [15:0] out_s903;
wire  [15:0] out_s904;
wire  [15:0] out_s905;
wire  [15:0] out_s906;
wire  [15:0] out_s907;
wire  [15:0] out_s908;
wire  [15:0] out_s909;
wire  [15:0] out_s910;
wire  [15:0] out_s911;
wire  [15:0] out_s912;
wire  [15:0] out_s913;
wire  [15:0] out_s914;
wire  [15:0] out_s915;
wire  [15:0] out_s916;
wire  [15:0] out_s917;
wire  [15:0] out_s918;
wire  [15:0] out_s919;
wire  [15:0] out_s920;
wire  [15:0] out_s921;
wire  [15:0] out_s922;
wire  [15:0] out_s923;
wire  [15:0] out_s924;
wire  [15:0] out_s925;
wire  [15:0] out_s926;
wire  [15:0] out_s927;
wire  [15:0] out_s928;
wire  [15:0] out_s929;
wire  [15:0] out_s930;
wire  [15:0] out_s931;
wire  [15:0] out_s932;
wire  [15:0] out_s933;
wire  [15:0] out_s934;
wire  [15:0] out_s935;
wire  [15:0] out_s936;
wire  [15:0] out_s937;
wire  [15:0] out_s938;
wire  [15:0] out_s939;
wire  [15:0] out_s940;
wire  [15:0] out_s941;
wire  [15:0] out_s942;
wire  [15:0] out_s943;
wire  [15:0] out_s944;
wire  [15:0] out_s945;
wire  [15:0] out_s946;
wire  [15:0] out_s947;
wire  [15:0] out_s948;
wire  [15:0] out_s949;
wire  [15:0] out_s950;
wire  [15:0] out_s951;
wire  [15:0] out_s952;
wire  [15:0] out_s953;
wire  [15:0] out_s954;
wire  [15:0] out_s955;
wire  [15:0] out_s956;
wire  [15:0] out_s957;
wire  [15:0] out_s958;
wire  [15:0] out_s959;
wire  [15:0] out_s960;
wire  [15:0] out_s961;
wire  [15:0] out_s962;
wire  [15:0] out_s963;
wire  [15:0] out_s964;
wire  [15:0] out_s965;
wire  [15:0] out_s966;
wire  [15:0] out_s967;
wire  [15:0] out_s968;
wire  [15:0] out_s969;
wire  [15:0] out_s970;
wire  [15:0] out_s971;
wire  [15:0] out_s972;
wire  [15:0] out_s973;
wire  [15:0] out_s974;
wire  [15:0] out_s975;
wire  [15:0] out_s976;
wire  [15:0] out_s977;
wire  [15:0] out_s978;
wire  [15:0] out_s979;
wire  [15:0] out_s980;
wire  [15:0] out_s981;
wire  [15:0] out_s982;
wire  [15:0] out_s983;
wire  [15:0] out_s984;
wire  [15:0] out_s985;
wire  [15:0] out_s986;
wire  [15:0] out_s987;
wire  [15:0] out_s988;
wire  [15:0] out_s989;
wire  [15:0] out_s990;
wire  [15:0] out_s991;
wire  [15:0] out_s992;
wire  [15:0] out_s993;
wire  [15:0] out_s994;
wire  [15:0] out_s995;
wire  [15:0] out_s996;
wire  [15:0] out_s997;
wire  [15:0] out_s998;
wire  [15:0] out_s999;
wire  [15:0] out_s1000;
wire  [15:0] out_s1001;
wire  [15:0] out_s1002;
wire  [15:0] out_s1003;
wire  [15:0] out_s1004;
wire  [15:0] out_s1005;
wire  [15:0] out_s1006;
wire  [15:0] out_s1007;
wire  [15:0] out_s1008;
wire  [15:0] out_s1009;
wire  [15:0] out_s1010;
wire  [15:0] out_s1011;
wire  [15:0] out_s1012;
wire  [15:0] out_s1013;
wire  [15:0] out_s1014;
wire  [15:0] out_s1015;
wire  [15:0] out_s1016;
wire  [15:0] out_s1017;
wire  [15:0] out_s1018;
wire  [15:0] out_s1019;
wire  [15:0] out_s1020;
wire  [15:0] out_s1021;
wire  [15:0] out_s1022;
wire  [15:0] out_s1023;

wire  [15:0] out_e0;
wire  [15:0] out_e1;
wire  [15:0] out_e2;
wire  [15:0] out_e3;
wire  [15:0] out_e4;
wire  [15:0] out_e5;
wire  [15:0] out_e6;
wire  [15:0] out_e7;
wire  [15:0] out_e8;
wire  [15:0] out_e9;
wire  [15:0] out_e10;
wire  [15:0] out_e11;
wire  [15:0] out_e12;
wire  [15:0] out_e13;
wire  [15:0] out_e14;
wire  [15:0] out_e15;
wire  [15:0] out_e16;
wire  [15:0] out_e17;
wire  [15:0] out_e18;
wire  [15:0] out_e19;
wire  [15:0] out_e20;
wire  [15:0] out_e21;
wire  [15:0] out_e22;
wire  [15:0] out_e23;
wire  [15:0] out_e24;
wire  [15:0] out_e25;
wire  [15:0] out_e26;
wire  [15:0] out_e27;
wire  [15:0] out_e28;
wire  [15:0] out_e29;
wire  [15:0] out_e30;
wire  [15:0] out_e31;
wire  [15:0] out_e32;
wire  [15:0] out_e33;
wire  [15:0] out_e34;
wire  [15:0] out_e35;
wire  [15:0] out_e36;
wire  [15:0] out_e37;
wire  [15:0] out_e38;
wire  [15:0] out_e39;
wire  [15:0] out_e40;
wire  [15:0] out_e41;
wire  [15:0] out_e42;
wire  [15:0] out_e43;
wire  [15:0] out_e44;
wire  [15:0] out_e45;
wire  [15:0] out_e46;
wire  [15:0] out_e47;
wire  [15:0] out_e48;
wire  [15:0] out_e49;
wire  [15:0] out_e50;
wire  [15:0] out_e51;
wire  [15:0] out_e52;
wire  [15:0] out_e53;
wire  [15:0] out_e54;
wire  [15:0] out_e55;
wire  [15:0] out_e56;
wire  [15:0] out_e57;
wire  [15:0] out_e58;
wire  [15:0] out_e59;
wire  [15:0] out_e60;
wire  [15:0] out_e61;
wire  [15:0] out_e62;
wire  [15:0] out_e63;
wire  [15:0] out_e64;
wire  [15:0] out_e65;
wire  [15:0] out_e66;
wire  [15:0] out_e67;
wire  [15:0] out_e68;
wire  [15:0] out_e69;
wire  [15:0] out_e70;
wire  [15:0] out_e71;
wire  [15:0] out_e72;
wire  [15:0] out_e73;
wire  [15:0] out_e74;
wire  [15:0] out_e75;
wire  [15:0] out_e76;
wire  [15:0] out_e77;
wire  [15:0] out_e78;
wire  [15:0] out_e79;
wire  [15:0] out_e80;
wire  [15:0] out_e81;
wire  [15:0] out_e82;
wire  [15:0] out_e83;
wire  [15:0] out_e84;
wire  [15:0] out_e85;
wire  [15:0] out_e86;
wire  [15:0] out_e87;
wire  [15:0] out_e88;
wire  [15:0] out_e89;
wire  [15:0] out_e90;
wire  [15:0] out_e91;
wire  [15:0] out_e92;
wire  [15:0] out_e93;
wire  [15:0] out_e94;
wire  [15:0] out_e95;
wire  [15:0] out_e96;
wire  [15:0] out_e97;
wire  [15:0] out_e98;
wire  [15:0] out_e99;
wire  [15:0] out_e100;
wire  [15:0] out_e101;
wire  [15:0] out_e102;
wire  [15:0] out_e103;
wire  [15:0] out_e104;
wire  [15:0] out_e105;
wire  [15:0] out_e106;
wire  [15:0] out_e107;
wire  [15:0] out_e108;
wire  [15:0] out_e109;
wire  [15:0] out_e110;
wire  [15:0] out_e111;
wire  [15:0] out_e112;
wire  [15:0] out_e113;
wire  [15:0] out_e114;
wire  [15:0] out_e115;
wire  [15:0] out_e116;
wire  [15:0] out_e117;
wire  [15:0] out_e118;
wire  [15:0] out_e119;
wire  [15:0] out_e120;
wire  [15:0] out_e121;
wire  [15:0] out_e122;
wire  [15:0] out_e123;
wire  [15:0] out_e124;
wire  [15:0] out_e125;
wire  [15:0] out_e126;
wire  [15:0] out_e127;
wire  [15:0] out_e128;
wire  [15:0] out_e129;
wire  [15:0] out_e130;
wire  [15:0] out_e131;
wire  [15:0] out_e132;
wire  [15:0] out_e133;
wire  [15:0] out_e134;
wire  [15:0] out_e135;
wire  [15:0] out_e136;
wire  [15:0] out_e137;
wire  [15:0] out_e138;
wire  [15:0] out_e139;
wire  [15:0] out_e140;
wire  [15:0] out_e141;
wire  [15:0] out_e142;
wire  [15:0] out_e143;
wire  [15:0] out_e144;
wire  [15:0] out_e145;
wire  [15:0] out_e146;
wire  [15:0] out_e147;
wire  [15:0] out_e148;
wire  [15:0] out_e149;
wire  [15:0] out_e150;
wire  [15:0] out_e151;
wire  [15:0] out_e152;
wire  [15:0] out_e153;
wire  [15:0] out_e154;
wire  [15:0] out_e155;
wire  [15:0] out_e156;
wire  [15:0] out_e157;
wire  [15:0] out_e158;
wire  [15:0] out_e159;
wire  [15:0] out_e160;
wire  [15:0] out_e161;
wire  [15:0] out_e162;
wire  [15:0] out_e163;
wire  [15:0] out_e164;
wire  [15:0] out_e165;
wire  [15:0] out_e166;
wire  [15:0] out_e167;
wire  [15:0] out_e168;
wire  [15:0] out_e169;
wire  [15:0] out_e170;
wire  [15:0] out_e171;
wire  [15:0] out_e172;
wire  [15:0] out_e173;
wire  [15:0] out_e174;
wire  [15:0] out_e175;
wire  [15:0] out_e176;
wire  [15:0] out_e177;
wire  [15:0] out_e178;
wire  [15:0] out_e179;
wire  [15:0] out_e180;
wire  [15:0] out_e181;
wire  [15:0] out_e182;
wire  [15:0] out_e183;
wire  [15:0] out_e184;
wire  [15:0] out_e185;
wire  [15:0] out_e186;
wire  [15:0] out_e187;
wire  [15:0] out_e188;
wire  [15:0] out_e189;
wire  [15:0] out_e190;
wire  [15:0] out_e191;
wire  [15:0] out_e192;
wire  [15:0] out_e193;
wire  [15:0] out_e194;
wire  [15:0] out_e195;
wire  [15:0] out_e196;
wire  [15:0] out_e197;
wire  [15:0] out_e198;
wire  [15:0] out_e199;
wire  [15:0] out_e200;
wire  [15:0] out_e201;
wire  [15:0] out_e202;
wire  [15:0] out_e203;
wire  [15:0] out_e204;
wire  [15:0] out_e205;
wire  [15:0] out_e206;
wire  [15:0] out_e207;
wire  [15:0] out_e208;
wire  [15:0] out_e209;
wire  [15:0] out_e210;
wire  [15:0] out_e211;
wire  [15:0] out_e212;
wire  [15:0] out_e213;
wire  [15:0] out_e214;
wire  [15:0] out_e215;
wire  [15:0] out_e216;
wire  [15:0] out_e217;
wire  [15:0] out_e218;
wire  [15:0] out_e219;
wire  [15:0] out_e220;
wire  [15:0] out_e221;
wire  [15:0] out_e222;
wire  [15:0] out_e223;
wire  [15:0] out_e224;
wire  [15:0] out_e225;
wire  [15:0] out_e226;
wire  [15:0] out_e227;
wire  [15:0] out_e228;
wire  [15:0] out_e229;
wire  [15:0] out_e230;
wire  [15:0] out_e231;
wire  [15:0] out_e232;
wire  [15:0] out_e233;
wire  [15:0] out_e234;
wire  [15:0] out_e235;
wire  [15:0] out_e236;
wire  [15:0] out_e237;
wire  [15:0] out_e238;
wire  [15:0] out_e239;
wire  [15:0] out_e240;
wire  [15:0] out_e241;
wire  [15:0] out_e242;
wire  [15:0] out_e243;
wire  [15:0] out_e244;
wire  [15:0] out_e245;
wire  [15:0] out_e246;
wire  [15:0] out_e247;
wire  [15:0] out_e248;
wire  [15:0] out_e249;
wire  [15:0] out_e250;
wire  [15:0] out_e251;
wire  [15:0] out_e252;
wire  [15:0] out_e253;
wire  [15:0] out_e254;
wire  [15:0] out_e255;
wire  [15:0] out_e256;
wire  [15:0] out_e257;
wire  [15:0] out_e258;
wire  [15:0] out_e259;
wire  [15:0] out_e260;
wire  [15:0] out_e261;
wire  [15:0] out_e262;
wire  [15:0] out_e263;
wire  [15:0] out_e264;
wire  [15:0] out_e265;
wire  [15:0] out_e266;
wire  [15:0] out_e267;
wire  [15:0] out_e268;
wire  [15:0] out_e269;
wire  [15:0] out_e270;
wire  [15:0] out_e271;
wire  [15:0] out_e272;
wire  [15:0] out_e273;
wire  [15:0] out_e274;
wire  [15:0] out_e275;
wire  [15:0] out_e276;
wire  [15:0] out_e277;
wire  [15:0] out_e278;
wire  [15:0] out_e279;
wire  [15:0] out_e280;
wire  [15:0] out_e281;
wire  [15:0] out_e282;
wire  [15:0] out_e283;
wire  [15:0] out_e284;
wire  [15:0] out_e285;
wire  [15:0] out_e286;
wire  [15:0] out_e287;
wire  [15:0] out_e288;
wire  [15:0] out_e289;
wire  [15:0] out_e290;
wire  [15:0] out_e291;
wire  [15:0] out_e292;
wire  [15:0] out_e293;
wire  [15:0] out_e294;
wire  [15:0] out_e295;
wire  [15:0] out_e296;
wire  [15:0] out_e297;
wire  [15:0] out_e298;
wire  [15:0] out_e299;
wire  [15:0] out_e300;
wire  [15:0] out_e301;
wire  [15:0] out_e302;
wire  [15:0] out_e303;
wire  [15:0] out_e304;
wire  [15:0] out_e305;
wire  [15:0] out_e306;
wire  [15:0] out_e307;
wire  [15:0] out_e308;
wire  [15:0] out_e309;
wire  [15:0] out_e310;
wire  [15:0] out_e311;
wire  [15:0] out_e312;
wire  [15:0] out_e313;
wire  [15:0] out_e314;
wire  [15:0] out_e315;
wire  [15:0] out_e316;
wire  [15:0] out_e317;
wire  [15:0] out_e318;
wire  [15:0] out_e319;
wire  [15:0] out_e320;
wire  [15:0] out_e321;
wire  [15:0] out_e322;
wire  [15:0] out_e323;
wire  [15:0] out_e324;
wire  [15:0] out_e325;
wire  [15:0] out_e326;
wire  [15:0] out_e327;
wire  [15:0] out_e328;
wire  [15:0] out_e329;
wire  [15:0] out_e330;
wire  [15:0] out_e331;
wire  [15:0] out_e332;
wire  [15:0] out_e333;
wire  [15:0] out_e334;
wire  [15:0] out_e335;
wire  [15:0] out_e336;
wire  [15:0] out_e337;
wire  [15:0] out_e338;
wire  [15:0] out_e339;
wire  [15:0] out_e340;
wire  [15:0] out_e341;
wire  [15:0] out_e342;
wire  [15:0] out_e343;
wire  [15:0] out_e344;
wire  [15:0] out_e345;
wire  [15:0] out_e346;
wire  [15:0] out_e347;
wire  [15:0] out_e348;
wire  [15:0] out_e349;
wire  [15:0] out_e350;
wire  [15:0] out_e351;
wire  [15:0] out_e352;
wire  [15:0] out_e353;
wire  [15:0] out_e354;
wire  [15:0] out_e355;
wire  [15:0] out_e356;
wire  [15:0] out_e357;
wire  [15:0] out_e358;
wire  [15:0] out_e359;
wire  [15:0] out_e360;
wire  [15:0] out_e361;
wire  [15:0] out_e362;
wire  [15:0] out_e363;
wire  [15:0] out_e364;
wire  [15:0] out_e365;
wire  [15:0] out_e366;
wire  [15:0] out_e367;
wire  [15:0] out_e368;
wire  [15:0] out_e369;
wire  [15:0] out_e370;
wire  [15:0] out_e371;
wire  [15:0] out_e372;
wire  [15:0] out_e373;
wire  [15:0] out_e374;
wire  [15:0] out_e375;
wire  [15:0] out_e376;
wire  [15:0] out_e377;
wire  [15:0] out_e378;
wire  [15:0] out_e379;
wire  [15:0] out_e380;
wire  [15:0] out_e381;
wire  [15:0] out_e382;
wire  [15:0] out_e383;
wire  [15:0] out_e384;
wire  [15:0] out_e385;
wire  [15:0] out_e386;
wire  [15:0] out_e387;
wire  [15:0] out_e388;
wire  [15:0] out_e389;
wire  [15:0] out_e390;
wire  [15:0] out_e391;
wire  [15:0] out_e392;
wire  [15:0] out_e393;
wire  [15:0] out_e394;
wire  [15:0] out_e395;
wire  [15:0] out_e396;
wire  [15:0] out_e397;
wire  [15:0] out_e398;
wire  [15:0] out_e399;
wire  [15:0] out_e400;
wire  [15:0] out_e401;
wire  [15:0] out_e402;
wire  [15:0] out_e403;
wire  [15:0] out_e404;
wire  [15:0] out_e405;
wire  [15:0] out_e406;
wire  [15:0] out_e407;
wire  [15:0] out_e408;
wire  [15:0] out_e409;
wire  [15:0] out_e410;
wire  [15:0] out_e411;
wire  [15:0] out_e412;
wire  [15:0] out_e413;
wire  [15:0] out_e414;
wire  [15:0] out_e415;
wire  [15:0] out_e416;
wire  [15:0] out_e417;
wire  [15:0] out_e418;
wire  [15:0] out_e419;
wire  [15:0] out_e420;
wire  [15:0] out_e421;
wire  [15:0] out_e422;
wire  [15:0] out_e423;
wire  [15:0] out_e424;
wire  [15:0] out_e425;
wire  [15:0] out_e426;
wire  [15:0] out_e427;
wire  [15:0] out_e428;
wire  [15:0] out_e429;
wire  [15:0] out_e430;
wire  [15:0] out_e431;
wire  [15:0] out_e432;
wire  [15:0] out_e433;
wire  [15:0] out_e434;
wire  [15:0] out_e435;
wire  [15:0] out_e436;
wire  [15:0] out_e437;
wire  [15:0] out_e438;
wire  [15:0] out_e439;
wire  [15:0] out_e440;
wire  [15:0] out_e441;
wire  [15:0] out_e442;
wire  [15:0] out_e443;
wire  [15:0] out_e444;
wire  [15:0] out_e445;
wire  [15:0] out_e446;
wire  [15:0] out_e447;
wire  [15:0] out_e448;
wire  [15:0] out_e449;
wire  [15:0] out_e450;
wire  [15:0] out_e451;
wire  [15:0] out_e452;
wire  [15:0] out_e453;
wire  [15:0] out_e454;
wire  [15:0] out_e455;
wire  [15:0] out_e456;
wire  [15:0] out_e457;
wire  [15:0] out_e458;
wire  [15:0] out_e459;
wire  [15:0] out_e460;
wire  [15:0] out_e461;
wire  [15:0] out_e462;
wire  [15:0] out_e463;
wire  [15:0] out_e464;
wire  [15:0] out_e465;
wire  [15:0] out_e466;
wire  [15:0] out_e467;
wire  [15:0] out_e468;
wire  [15:0] out_e469;
wire  [15:0] out_e470;
wire  [15:0] out_e471;
wire  [15:0] out_e472;
wire  [15:0] out_e473;
wire  [15:0] out_e474;
wire  [15:0] out_e475;
wire  [15:0] out_e476;
wire  [15:0] out_e477;
wire  [15:0] out_e478;
wire  [15:0] out_e479;
wire  [15:0] out_e480;
wire  [15:0] out_e481;
wire  [15:0] out_e482;
wire  [15:0] out_e483;
wire  [15:0] out_e484;
wire  [15:0] out_e485;
wire  [15:0] out_e486;
wire  [15:0] out_e487;
wire  [15:0] out_e488;
wire  [15:0] out_e489;
wire  [15:0] out_e490;
wire  [15:0] out_e491;
wire  [15:0] out_e492;
wire  [15:0] out_e493;
wire  [15:0] out_e494;
wire  [15:0] out_e495;
wire  [15:0] out_e496;
wire  [15:0] out_e497;
wire  [15:0] out_e498;
wire  [15:0] out_e499;
wire  [15:0] out_e500;
wire  [15:0] out_e501;
wire  [15:0] out_e502;
wire  [15:0] out_e503;
wire  [15:0] out_e504;
wire  [15:0] out_e505;
wire  [15:0] out_e506;
wire  [15:0] out_e507;
wire  [15:0] out_e508;
wire  [15:0] out_e509;
wire  [15:0] out_e510;
wire  [15:0] out_e511;
wire  [15:0] out_e512;
wire  [15:0] out_e513;
wire  [15:0] out_e514;
wire  [15:0] out_e515;
wire  [15:0] out_e516;
wire  [15:0] out_e517;
wire  [15:0] out_e518;
wire  [15:0] out_e519;
wire  [15:0] out_e520;
wire  [15:0] out_e521;
wire  [15:0] out_e522;
wire  [15:0] out_e523;
wire  [15:0] out_e524;
wire  [15:0] out_e525;
wire  [15:0] out_e526;
wire  [15:0] out_e527;
wire  [15:0] out_e528;
wire  [15:0] out_e529;
wire  [15:0] out_e530;
wire  [15:0] out_e531;
wire  [15:0] out_e532;
wire  [15:0] out_e533;
wire  [15:0] out_e534;
wire  [15:0] out_e535;
wire  [15:0] out_e536;
wire  [15:0] out_e537;
wire  [15:0] out_e538;
wire  [15:0] out_e539;
wire  [15:0] out_e540;
wire  [15:0] out_e541;
wire  [15:0] out_e542;
wire  [15:0] out_e543;
wire  [15:0] out_e544;
wire  [15:0] out_e545;
wire  [15:0] out_e546;
wire  [15:0] out_e547;
wire  [15:0] out_e548;
wire  [15:0] out_e549;
wire  [15:0] out_e550;
wire  [15:0] out_e551;
wire  [15:0] out_e552;
wire  [15:0] out_e553;
wire  [15:0] out_e554;
wire  [15:0] out_e555;
wire  [15:0] out_e556;
wire  [15:0] out_e557;
wire  [15:0] out_e558;
wire  [15:0] out_e559;
wire  [15:0] out_e560;
wire  [15:0] out_e561;
wire  [15:0] out_e562;
wire  [15:0] out_e563;
wire  [15:0] out_e564;
wire  [15:0] out_e565;
wire  [15:0] out_e566;
wire  [15:0] out_e567;
wire  [15:0] out_e568;
wire  [15:0] out_e569;
wire  [15:0] out_e570;
wire  [15:0] out_e571;
wire  [15:0] out_e572;
wire  [15:0] out_e573;
wire  [15:0] out_e574;
wire  [15:0] out_e575;
wire  [15:0] out_e576;
wire  [15:0] out_e577;
wire  [15:0] out_e578;
wire  [15:0] out_e579;
wire  [15:0] out_e580;
wire  [15:0] out_e581;
wire  [15:0] out_e582;
wire  [15:0] out_e583;
wire  [15:0] out_e584;
wire  [15:0] out_e585;
wire  [15:0] out_e586;
wire  [15:0] out_e587;
wire  [15:0] out_e588;
wire  [15:0] out_e589;
wire  [15:0] out_e590;
wire  [15:0] out_e591;
wire  [15:0] out_e592;
wire  [15:0] out_e593;
wire  [15:0] out_e594;
wire  [15:0] out_e595;
wire  [15:0] out_e596;
wire  [15:0] out_e597;
wire  [15:0] out_e598;
wire  [15:0] out_e599;
wire  [15:0] out_e600;
wire  [15:0] out_e601;
wire  [15:0] out_e602;
wire  [15:0] out_e603;
wire  [15:0] out_e604;
wire  [15:0] out_e605;
wire  [15:0] out_e606;
wire  [15:0] out_e607;
wire  [15:0] out_e608;
wire  [15:0] out_e609;
wire  [15:0] out_e610;
wire  [15:0] out_e611;
wire  [15:0] out_e612;
wire  [15:0] out_e613;
wire  [15:0] out_e614;
wire  [15:0] out_e615;
wire  [15:0] out_e616;
wire  [15:0] out_e617;
wire  [15:0] out_e618;
wire  [15:0] out_e619;
wire  [15:0] out_e620;
wire  [15:0] out_e621;
wire  [15:0] out_e622;
wire  [15:0] out_e623;
wire  [15:0] out_e624;
wire  [15:0] out_e625;
wire  [15:0] out_e626;
wire  [15:0] out_e627;
wire  [15:0] out_e628;
wire  [15:0] out_e629;
wire  [15:0] out_e630;
wire  [15:0] out_e631;
wire  [15:0] out_e632;
wire  [15:0] out_e633;
wire  [15:0] out_e634;
wire  [15:0] out_e635;
wire  [15:0] out_e636;
wire  [15:0] out_e637;
wire  [15:0] out_e638;
wire  [15:0] out_e639;
wire  [15:0] out_e640;
wire  [15:0] out_e641;
wire  [15:0] out_e642;
wire  [15:0] out_e643;
wire  [15:0] out_e644;
wire  [15:0] out_e645;
wire  [15:0] out_e646;
wire  [15:0] out_e647;
wire  [15:0] out_e648;
wire  [15:0] out_e649;
wire  [15:0] out_e650;
wire  [15:0] out_e651;
wire  [15:0] out_e652;
wire  [15:0] out_e653;
wire  [15:0] out_e654;
wire  [15:0] out_e655;
wire  [15:0] out_e656;
wire  [15:0] out_e657;
wire  [15:0] out_e658;
wire  [15:0] out_e659;
wire  [15:0] out_e660;
wire  [15:0] out_e661;
wire  [15:0] out_e662;
wire  [15:0] out_e663;
wire  [15:0] out_e664;
wire  [15:0] out_e665;
wire  [15:0] out_e666;
wire  [15:0] out_e667;
wire  [15:0] out_e668;
wire  [15:0] out_e669;
wire  [15:0] out_e670;
wire  [15:0] out_e671;
wire  [15:0] out_e672;
wire  [15:0] out_e673;
wire  [15:0] out_e674;
wire  [15:0] out_e675;
wire  [15:0] out_e676;
wire  [15:0] out_e677;
wire  [15:0] out_e678;
wire  [15:0] out_e679;
wire  [15:0] out_e680;
wire  [15:0] out_e681;
wire  [15:0] out_e682;
wire  [15:0] out_e683;
wire  [15:0] out_e684;
wire  [15:0] out_e685;
wire  [15:0] out_e686;
wire  [15:0] out_e687;
wire  [15:0] out_e688;
wire  [15:0] out_e689;
wire  [15:0] out_e690;
wire  [15:0] out_e691;
wire  [15:0] out_e692;
wire  [15:0] out_e693;
wire  [15:0] out_e694;
wire  [15:0] out_e695;
wire  [15:0] out_e696;
wire  [15:0] out_e697;
wire  [15:0] out_e698;
wire  [15:0] out_e699;
wire  [15:0] out_e700;
wire  [15:0] out_e701;
wire  [15:0] out_e702;
wire  [15:0] out_e703;
wire  [15:0] out_e704;
wire  [15:0] out_e705;
wire  [15:0] out_e706;
wire  [15:0] out_e707;
wire  [15:0] out_e708;
wire  [15:0] out_e709;
wire  [15:0] out_e710;
wire  [15:0] out_e711;
wire  [15:0] out_e712;
wire  [15:0] out_e713;
wire  [15:0] out_e714;
wire  [15:0] out_e715;
wire  [15:0] out_e716;
wire  [15:0] out_e717;
wire  [15:0] out_e718;
wire  [15:0] out_e719;
wire  [15:0] out_e720;
wire  [15:0] out_e721;
wire  [15:0] out_e722;
wire  [15:0] out_e723;
wire  [15:0] out_e724;
wire  [15:0] out_e725;
wire  [15:0] out_e726;
wire  [15:0] out_e727;
wire  [15:0] out_e728;
wire  [15:0] out_e729;
wire  [15:0] out_e730;
wire  [15:0] out_e731;
wire  [15:0] out_e732;
wire  [15:0] out_e733;
wire  [15:0] out_e734;
wire  [15:0] out_e735;
wire  [15:0] out_e736;
wire  [15:0] out_e737;
wire  [15:0] out_e738;
wire  [15:0] out_e739;
wire  [15:0] out_e740;
wire  [15:0] out_e741;
wire  [15:0] out_e742;
wire  [15:0] out_e743;
wire  [15:0] out_e744;
wire  [15:0] out_e745;
wire  [15:0] out_e746;
wire  [15:0] out_e747;
wire  [15:0] out_e748;
wire  [15:0] out_e749;
wire  [15:0] out_e750;
wire  [15:0] out_e751;
wire  [15:0] out_e752;
wire  [15:0] out_e753;
wire  [15:0] out_e754;
wire  [15:0] out_e755;
wire  [15:0] out_e756;
wire  [15:0] out_e757;
wire  [15:0] out_e758;
wire  [15:0] out_e759;
wire  [15:0] out_e760;
wire  [15:0] out_e761;
wire  [15:0] out_e762;
wire  [15:0] out_e763;
wire  [15:0] out_e764;
wire  [15:0] out_e765;
wire  [15:0] out_e766;
wire  [15:0] out_e767;
wire  [15:0] out_e768;
wire  [15:0] out_e769;
wire  [15:0] out_e770;
wire  [15:0] out_e771;
wire  [15:0] out_e772;
wire  [15:0] out_e773;
wire  [15:0] out_e774;
wire  [15:0] out_e775;
wire  [15:0] out_e776;
wire  [15:0] out_e777;
wire  [15:0] out_e778;
wire  [15:0] out_e779;
wire  [15:0] out_e780;
wire  [15:0] out_e781;
wire  [15:0] out_e782;
wire  [15:0] out_e783;
wire  [15:0] out_e784;
wire  [15:0] out_e785;
wire  [15:0] out_e786;
wire  [15:0] out_e787;
wire  [15:0] out_e788;
wire  [15:0] out_e789;
wire  [15:0] out_e790;
wire  [15:0] out_e791;
wire  [15:0] out_e792;
wire  [15:0] out_e793;
wire  [15:0] out_e794;
wire  [15:0] out_e795;
wire  [15:0] out_e796;
wire  [15:0] out_e797;
wire  [15:0] out_e798;
wire  [15:0] out_e799;
wire  [15:0] out_e800;
wire  [15:0] out_e801;
wire  [15:0] out_e802;
wire  [15:0] out_e803;
wire  [15:0] out_e804;
wire  [15:0] out_e805;
wire  [15:0] out_e806;
wire  [15:0] out_e807;
wire  [15:0] out_e808;
wire  [15:0] out_e809;
wire  [15:0] out_e810;
wire  [15:0] out_e811;
wire  [15:0] out_e812;
wire  [15:0] out_e813;
wire  [15:0] out_e814;
wire  [15:0] out_e815;
wire  [15:0] out_e816;
wire  [15:0] out_e817;
wire  [15:0] out_e818;
wire  [15:0] out_e819;
wire  [15:0] out_e820;
wire  [15:0] out_e821;
wire  [15:0] out_e822;
wire  [15:0] out_e823;
wire  [15:0] out_e824;
wire  [15:0] out_e825;
wire  [15:0] out_e826;
wire  [15:0] out_e827;
wire  [15:0] out_e828;
wire  [15:0] out_e829;
wire  [15:0] out_e830;
wire  [15:0] out_e831;
wire  [15:0] out_e832;
wire  [15:0] out_e833;
wire  [15:0] out_e834;
wire  [15:0] out_e835;
wire  [15:0] out_e836;
wire  [15:0] out_e837;
wire  [15:0] out_e838;
wire  [15:0] out_e839;
wire  [15:0] out_e840;
wire  [15:0] out_e841;
wire  [15:0] out_e842;
wire  [15:0] out_e843;
wire  [15:0] out_e844;
wire  [15:0] out_e845;
wire  [15:0] out_e846;
wire  [15:0] out_e847;
wire  [15:0] out_e848;
wire  [15:0] out_e849;
wire  [15:0] out_e850;
wire  [15:0] out_e851;
wire  [15:0] out_e852;
wire  [15:0] out_e853;
wire  [15:0] out_e854;
wire  [15:0] out_e855;
wire  [15:0] out_e856;
wire  [15:0] out_e857;
wire  [15:0] out_e858;
wire  [15:0] out_e859;
wire  [15:0] out_e860;
wire  [15:0] out_e861;
wire  [15:0] out_e862;
wire  [15:0] out_e863;
wire  [15:0] out_e864;
wire  [15:0] out_e865;
wire  [15:0] out_e866;
wire  [15:0] out_e867;
wire  [15:0] out_e868;
wire  [15:0] out_e869;
wire  [15:0] out_e870;
wire  [15:0] out_e871;
wire  [15:0] out_e872;
wire  [15:0] out_e873;
wire  [15:0] out_e874;
wire  [15:0] out_e875;
wire  [15:0] out_e876;
wire  [15:0] out_e877;
wire  [15:0] out_e878;
wire  [15:0] out_e879;
wire  [15:0] out_e880;
wire  [15:0] out_e881;
wire  [15:0] out_e882;
wire  [15:0] out_e883;
wire  [15:0] out_e884;
wire  [15:0] out_e885;
wire  [15:0] out_e886;
wire  [15:0] out_e887;
wire  [15:0] out_e888;
wire  [15:0] out_e889;
wire  [15:0] out_e890;
wire  [15:0] out_e891;
wire  [15:0] out_e892;
wire  [15:0] out_e893;
wire  [15:0] out_e894;
wire  [15:0] out_e895;
wire  [15:0] out_e896;
wire  [15:0] out_e897;
wire  [15:0] out_e898;
wire  [15:0] out_e899;
wire  [15:0] out_e900;
wire  [15:0] out_e901;
wire  [15:0] out_e902;
wire  [15:0] out_e903;
wire  [15:0] out_e904;
wire  [15:0] out_e905;
wire  [15:0] out_e906;
wire  [15:0] out_e907;
wire  [15:0] out_e908;
wire  [15:0] out_e909;
wire  [15:0] out_e910;
wire  [15:0] out_e911;
wire  [15:0] out_e912;
wire  [15:0] out_e913;
wire  [15:0] out_e914;
wire  [15:0] out_e915;
wire  [15:0] out_e916;
wire  [15:0] out_e917;
wire  [15:0] out_e918;
wire  [15:0] out_e919;
wire  [15:0] out_e920;
wire  [15:0] out_e921;
wire  [15:0] out_e922;
wire  [15:0] out_e923;
wire  [15:0] out_e924;
wire  [15:0] out_e925;
wire  [15:0] out_e926;
wire  [15:0] out_e927;
wire  [15:0] out_e928;
wire  [15:0] out_e929;
wire  [15:0] out_e930;
wire  [15:0] out_e931;
wire  [15:0] out_e932;
wire  [15:0] out_e933;
wire  [15:0] out_e934;
wire  [15:0] out_e935;
wire  [15:0] out_e936;
wire  [15:0] out_e937;
wire  [15:0] out_e938;
wire  [15:0] out_e939;
wire  [15:0] out_e940;
wire  [15:0] out_e941;
wire  [15:0] out_e942;
wire  [15:0] out_e943;
wire  [15:0] out_e944;
wire  [15:0] out_e945;
wire  [15:0] out_e946;
wire  [15:0] out_e947;
wire  [15:0] out_e948;
wire  [15:0] out_e949;
wire  [15:0] out_e950;
wire  [15:0] out_e951;
wire  [15:0] out_e952;
wire  [15:0] out_e953;
wire  [15:0] out_e954;
wire  [15:0] out_e955;
wire  [15:0] out_e956;
wire  [15:0] out_e957;
wire  [15:0] out_e958;
wire  [15:0] out_e959;
wire  [15:0] out_e960;
wire  [15:0] out_e961;
wire  [15:0] out_e962;
wire  [15:0] out_e963;
wire  [15:0] out_e964;
wire  [15:0] out_e965;
wire  [15:0] out_e966;
wire  [15:0] out_e967;
wire  [15:0] out_e968;
wire  [15:0] out_e969;
wire  [15:0] out_e970;
wire  [15:0] out_e971;
wire  [15:0] out_e972;
wire  [15:0] out_e973;
wire  [15:0] out_e974;
wire  [15:0] out_e975;
wire  [15:0] out_e976;
wire  [15:0] out_e977;
wire  [15:0] out_e978;
wire  [15:0] out_e979;
wire  [15:0] out_e980;
wire  [15:0] out_e981;
wire  [15:0] out_e982;
wire  [15:0] out_e983;
wire  [15:0] out_e984;
wire  [15:0] out_e985;
wire  [15:0] out_e986;
wire  [15:0] out_e987;
wire  [15:0] out_e988;
wire  [15:0] out_e989;
wire  [15:0] out_e990;
wire  [15:0] out_e991;
wire  [15:0] out_e992;
wire  [15:0] out_e993;
wire  [15:0] out_e994;
wire  [15:0] out_e995;
wire  [15:0] out_e996;
wire  [15:0] out_e997;
wire  [15:0] out_e998;
wire  [15:0] out_e999;
wire  [15:0] out_e1000;
wire  [15:0] out_e1001;
wire  [15:0] out_e1002;
wire  [15:0] out_e1003;
wire  [15:0] out_e1004;
wire  [15:0] out_e1005;
wire  [15:0] out_e1006;
wire  [15:0] out_e1007;
wire  [15:0] out_e1008;
wire  [15:0] out_e1009;
wire  [15:0] out_e1010;
wire  [15:0] out_e1011;
wire  [15:0] out_e1012;
wire  [15:0] out_e1013;
wire  [15:0] out_e1014;
wire  [15:0] out_e1015;
wire  [15:0] out_e1016;
wire  [15:0] out_e1017;
wire  [15:0] out_e1018;
wire  [15:0] out_e1019;
wire  [15:0] out_e1020;
wire  [15:0] out_e1021;
wire  [15:0] out_e1022;
wire  [15:0] out_e1023;

wire  [15:0] result0;
wire  [15:0] result1;
wire  [15:0] result2;
wire  [15:0] result3;
wire  [15:0] result4;
wire  [15:0] result5;
wire  [15:0] result6;
wire  [15:0] result7;
wire  [15:0] result8;
wire  [15:0] result9;
wire  [15:0] result10;
wire  [15:0] result11;
wire  [15:0] result12;
wire  [15:0] result13;
wire  [15:0] result14;
wire  [15:0] result15;
wire  [15:0] result16;
wire  [15:0] result17;
wire  [15:0] result18;
wire  [15:0] result19;
wire  [15:0] result20;
wire  [15:0] result21;
wire  [15:0] result22;
wire  [15:0] result23;
wire  [15:0] result24;
wire  [15:0] result25;
wire  [15:0] result26;
wire  [15:0] result27;
wire  [15:0] result28;
wire  [15:0] result29;
wire  [15:0] result30;
wire  [15:0] result31;
wire  [15:0] result32;
wire  [15:0] result33;
wire  [15:0] result34;
wire  [15:0] result35;
wire  [15:0] result36;
wire  [15:0] result37;
wire  [15:0] result38;
wire  [15:0] result39;
wire  [15:0] result40;
wire  [15:0] result41;
wire  [15:0] result42;
wire  [15:0] result43;
wire  [15:0] result44;
wire  [15:0] result45;
wire  [15:0] result46;
wire  [15:0] result47;
wire  [15:0] result48;
wire  [15:0] result49;
wire  [15:0] result50;
wire  [15:0] result51;
wire  [15:0] result52;
wire  [15:0] result53;
wire  [15:0] result54;
wire  [15:0] result55;
wire  [15:0] result56;
wire  [15:0] result57;
wire  [15:0] result58;
wire  [15:0] result59;
wire  [15:0] result60;
wire  [15:0] result61;
wire  [15:0] result62;
wire  [15:0] result63;
wire  [15:0] result64;
wire  [15:0] result65;
wire  [15:0] result66;
wire  [15:0] result67;
wire  [15:0] result68;
wire  [15:0] result69;
wire  [15:0] result70;
wire  [15:0] result71;
wire  [15:0] result72;
wire  [15:0] result73;
wire  [15:0] result74;
wire  [15:0] result75;
wire  [15:0] result76;
wire  [15:0] result77;
wire  [15:0] result78;
wire  [15:0] result79;
wire  [15:0] result80;
wire  [15:0] result81;
wire  [15:0] result82;
wire  [15:0] result83;
wire  [15:0] result84;
wire  [15:0] result85;
wire  [15:0] result86;
wire  [15:0] result87;
wire  [15:0] result88;
wire  [15:0] result89;
wire  [15:0] result90;
wire  [15:0] result91;
wire  [15:0] result92;
wire  [15:0] result93;
wire  [15:0] result94;
wire  [15:0] result95;
wire  [15:0] result96;
wire  [15:0] result97;
wire  [15:0] result98;
wire  [15:0] result99;
wire  [15:0] result100;
wire  [15:0] result101;
wire  [15:0] result102;
wire  [15:0] result103;
wire  [15:0] result104;
wire  [15:0] result105;
wire  [15:0] result106;
wire  [15:0] result107;
wire  [15:0] result108;
wire  [15:0] result109;
wire  [15:0] result110;
wire  [15:0] result111;
wire  [15:0] result112;
wire  [15:0] result113;
wire  [15:0] result114;
wire  [15:0] result115;
wire  [15:0] result116;
wire  [15:0] result117;
wire  [15:0] result118;
wire  [15:0] result119;
wire  [15:0] result120;
wire  [15:0] result121;
wire  [15:0] result122;
wire  [15:0] result123;
wire  [15:0] result124;
wire  [15:0] result125;
wire  [15:0] result126;
wire  [15:0] result127;
wire  [15:0] result128;
wire  [15:0] result129;
wire  [15:0] result130;
wire  [15:0] result131;
wire  [15:0] result132;
wire  [15:0] result133;
wire  [15:0] result134;
wire  [15:0] result135;
wire  [15:0] result136;
wire  [15:0] result137;
wire  [15:0] result138;
wire  [15:0] result139;
wire  [15:0] result140;
wire  [15:0] result141;
wire  [15:0] result142;
wire  [15:0] result143;
wire  [15:0] result144;
wire  [15:0] result145;
wire  [15:0] result146;
wire  [15:0] result147;
wire  [15:0] result148;
wire  [15:0] result149;
wire  [15:0] result150;
wire  [15:0] result151;
wire  [15:0] result152;
wire  [15:0] result153;
wire  [15:0] result154;
wire  [15:0] result155;
wire  [15:0] result156;
wire  [15:0] result157;
wire  [15:0] result158;
wire  [15:0] result159;
wire  [15:0] result160;
wire  [15:0] result161;
wire  [15:0] result162;
wire  [15:0] result163;
wire  [15:0] result164;
wire  [15:0] result165;
wire  [15:0] result166;
wire  [15:0] result167;
wire  [15:0] result168;
wire  [15:0] result169;
wire  [15:0] result170;
wire  [15:0] result171;
wire  [15:0] result172;
wire  [15:0] result173;
wire  [15:0] result174;
wire  [15:0] result175;
wire  [15:0] result176;
wire  [15:0] result177;
wire  [15:0] result178;
wire  [15:0] result179;
wire  [15:0] result180;
wire  [15:0] result181;
wire  [15:0] result182;
wire  [15:0] result183;
wire  [15:0] result184;
wire  [15:0] result185;
wire  [15:0] result186;
wire  [15:0] result187;
wire  [15:0] result188;
wire  [15:0] result189;
wire  [15:0] result190;
wire  [15:0] result191;
wire  [15:0] result192;
wire  [15:0] result193;
wire  [15:0] result194;
wire  [15:0] result195;
wire  [15:0] result196;
wire  [15:0] result197;
wire  [15:0] result198;
wire  [15:0] result199;
wire  [15:0] result200;
wire  [15:0] result201;
wire  [15:0] result202;
wire  [15:0] result203;
wire  [15:0] result204;
wire  [15:0] result205;
wire  [15:0] result206;
wire  [15:0] result207;
wire  [15:0] result208;
wire  [15:0] result209;
wire  [15:0] result210;
wire  [15:0] result211;
wire  [15:0] result212;
wire  [15:0] result213;
wire  [15:0] result214;
wire  [15:0] result215;
wire  [15:0] result216;
wire  [15:0] result217;
wire  [15:0] result218;
wire  [15:0] result219;
wire  [15:0] result220;
wire  [15:0] result221;
wire  [15:0] result222;
wire  [15:0] result223;
wire  [15:0] result224;
wire  [15:0] result225;
wire  [15:0] result226;
wire  [15:0] result227;
wire  [15:0] result228;
wire  [15:0] result229;
wire  [15:0] result230;
wire  [15:0] result231;
wire  [15:0] result232;
wire  [15:0] result233;
wire  [15:0] result234;
wire  [15:0] result235;
wire  [15:0] result236;
wire  [15:0] result237;
wire  [15:0] result238;
wire  [15:0] result239;
wire  [15:0] result240;
wire  [15:0] result241;
wire  [15:0] result242;
wire  [15:0] result243;
wire  [15:0] result244;
wire  [15:0] result245;
wire  [15:0] result246;
wire  [15:0] result247;
wire  [15:0] result248;
wire  [15:0] result249;
wire  [15:0] result250;
wire  [15:0] result251;
wire  [15:0] result252;
wire  [15:0] result253;
wire  [15:0] result254;
wire  [15:0] result255;
wire  [15:0] result256;
wire  [15:0] result257;
wire  [15:0] result258;
wire  [15:0] result259;
wire  [15:0] result260;
wire  [15:0] result261;
wire  [15:0] result262;
wire  [15:0] result263;
wire  [15:0] result264;
wire  [15:0] result265;
wire  [15:0] result266;
wire  [15:0] result267;
wire  [15:0] result268;
wire  [15:0] result269;
wire  [15:0] result270;
wire  [15:0] result271;
wire  [15:0] result272;
wire  [15:0] result273;
wire  [15:0] result274;
wire  [15:0] result275;
wire  [15:0] result276;
wire  [15:0] result277;
wire  [15:0] result278;
wire  [15:0] result279;
wire  [15:0] result280;
wire  [15:0] result281;
wire  [15:0] result282;
wire  [15:0] result283;
wire  [15:0] result284;
wire  [15:0] result285;
wire  [15:0] result286;
wire  [15:0] result287;
wire  [15:0] result288;
wire  [15:0] result289;
wire  [15:0] result290;
wire  [15:0] result291;
wire  [15:0] result292;
wire  [15:0] result293;
wire  [15:0] result294;
wire  [15:0] result295;
wire  [15:0] result296;
wire  [15:0] result297;
wire  [15:0] result298;
wire  [15:0] result299;
wire  [15:0] result300;
wire  [15:0] result301;
wire  [15:0] result302;
wire  [15:0] result303;
wire  [15:0] result304;
wire  [15:0] result305;
wire  [15:0] result306;
wire  [15:0] result307;
wire  [15:0] result308;
wire  [15:0] result309;
wire  [15:0] result310;
wire  [15:0] result311;
wire  [15:0] result312;
wire  [15:0] result313;
wire  [15:0] result314;
wire  [15:0] result315;
wire  [15:0] result316;
wire  [15:0] result317;
wire  [15:0] result318;
wire  [15:0] result319;
wire  [15:0] result320;
wire  [15:0] result321;
wire  [15:0] result322;
wire  [15:0] result323;
wire  [15:0] result324;
wire  [15:0] result325;
wire  [15:0] result326;
wire  [15:0] result327;
wire  [15:0] result328;
wire  [15:0] result329;
wire  [15:0] result330;
wire  [15:0] result331;
wire  [15:0] result332;
wire  [15:0] result333;
wire  [15:0] result334;
wire  [15:0] result335;
wire  [15:0] result336;
wire  [15:0] result337;
wire  [15:0] result338;
wire  [15:0] result339;
wire  [15:0] result340;
wire  [15:0] result341;
wire  [15:0] result342;
wire  [15:0] result343;
wire  [15:0] result344;
wire  [15:0] result345;
wire  [15:0] result346;
wire  [15:0] result347;
wire  [15:0] result348;
wire  [15:0] result349;
wire  [15:0] result350;
wire  [15:0] result351;
wire  [15:0] result352;
wire  [15:0] result353;
wire  [15:0] result354;
wire  [15:0] result355;
wire  [15:0] result356;
wire  [15:0] result357;
wire  [15:0] result358;
wire  [15:0] result359;
wire  [15:0] result360;
wire  [15:0] result361;
wire  [15:0] result362;
wire  [15:0] result363;
wire  [15:0] result364;
wire  [15:0] result365;
wire  [15:0] result366;
wire  [15:0] result367;
wire  [15:0] result368;
wire  [15:0] result369;
wire  [15:0] result370;
wire  [15:0] result371;
wire  [15:0] result372;
wire  [15:0] result373;
wire  [15:0] result374;
wire  [15:0] result375;
wire  [15:0] result376;
wire  [15:0] result377;
wire  [15:0] result378;
wire  [15:0] result379;
wire  [15:0] result380;
wire  [15:0] result381;
wire  [15:0] result382;
wire  [15:0] result383;
wire  [15:0] result384;
wire  [15:0] result385;
wire  [15:0] result386;
wire  [15:0] result387;
wire  [15:0] result388;
wire  [15:0] result389;
wire  [15:0] result390;
wire  [15:0] result391;
wire  [15:0] result392;
wire  [15:0] result393;
wire  [15:0] result394;
wire  [15:0] result395;
wire  [15:0] result396;
wire  [15:0] result397;
wire  [15:0] result398;
wire  [15:0] result399;
wire  [15:0] result400;
wire  [15:0] result401;
wire  [15:0] result402;
wire  [15:0] result403;
wire  [15:0] result404;
wire  [15:0] result405;
wire  [15:0] result406;
wire  [15:0] result407;
wire  [15:0] result408;
wire  [15:0] result409;
wire  [15:0] result410;
wire  [15:0] result411;
wire  [15:0] result412;
wire  [15:0] result413;
wire  [15:0] result414;
wire  [15:0] result415;
wire  [15:0] result416;
wire  [15:0] result417;
wire  [15:0] result418;
wire  [15:0] result419;
wire  [15:0] result420;
wire  [15:0] result421;
wire  [15:0] result422;
wire  [15:0] result423;
wire  [15:0] result424;
wire  [15:0] result425;
wire  [15:0] result426;
wire  [15:0] result427;
wire  [15:0] result428;
wire  [15:0] result429;
wire  [15:0] result430;
wire  [15:0] result431;
wire  [15:0] result432;
wire  [15:0] result433;
wire  [15:0] result434;
wire  [15:0] result435;
wire  [15:0] result436;
wire  [15:0] result437;
wire  [15:0] result438;
wire  [15:0] result439;
wire  [15:0] result440;
wire  [15:0] result441;
wire  [15:0] result442;
wire  [15:0] result443;
wire  [15:0] result444;
wire  [15:0] result445;
wire  [15:0] result446;
wire  [15:0] result447;
wire  [15:0] result448;
wire  [15:0] result449;
wire  [15:0] result450;
wire  [15:0] result451;
wire  [15:0] result452;
wire  [15:0] result453;
wire  [15:0] result454;
wire  [15:0] result455;
wire  [15:0] result456;
wire  [15:0] result457;
wire  [15:0] result458;
wire  [15:0] result459;
wire  [15:0] result460;
wire  [15:0] result461;
wire  [15:0] result462;
wire  [15:0] result463;
wire  [15:0] result464;
wire  [15:0] result465;
wire  [15:0] result466;
wire  [15:0] result467;
wire  [15:0] result468;
wire  [15:0] result469;
wire  [15:0] result470;
wire  [15:0] result471;
wire  [15:0] result472;
wire  [15:0] result473;
wire  [15:0] result474;
wire  [15:0] result475;
wire  [15:0] result476;
wire  [15:0] result477;
wire  [15:0] result478;
wire  [15:0] result479;
wire  [15:0] result480;
wire  [15:0] result481;
wire  [15:0] result482;
wire  [15:0] result483;
wire  [15:0] result484;
wire  [15:0] result485;
wire  [15:0] result486;
wire  [15:0] result487;
wire  [15:0] result488;
wire  [15:0] result489;
wire  [15:0] result490;
wire  [15:0] result491;
wire  [15:0] result492;
wire  [15:0] result493;
wire  [15:0] result494;
wire  [15:0] result495;
wire  [15:0] result496;
wire  [15:0] result497;
wire  [15:0] result498;
wire  [15:0] result499;
wire  [15:0] result500;
wire  [15:0] result501;
wire  [15:0] result502;
wire  [15:0] result503;
wire  [15:0] result504;
wire  [15:0] result505;
wire  [15:0] result506;
wire  [15:0] result507;
wire  [15:0] result508;
wire  [15:0] result509;
wire  [15:0] result510;
wire  [15:0] result511;
wire  [15:0] result512;
wire  [15:0] result513;
wire  [15:0] result514;
wire  [15:0] result515;
wire  [15:0] result516;
wire  [15:0] result517;
wire  [15:0] result518;
wire  [15:0] result519;
wire  [15:0] result520;
wire  [15:0] result521;
wire  [15:0] result522;
wire  [15:0] result523;
wire  [15:0] result524;
wire  [15:0] result525;
wire  [15:0] result526;
wire  [15:0] result527;
wire  [15:0] result528;
wire  [15:0] result529;
wire  [15:0] result530;
wire  [15:0] result531;
wire  [15:0] result532;
wire  [15:0] result533;
wire  [15:0] result534;
wire  [15:0] result535;
wire  [15:0] result536;
wire  [15:0] result537;
wire  [15:0] result538;
wire  [15:0] result539;
wire  [15:0] result540;
wire  [15:0] result541;
wire  [15:0] result542;
wire  [15:0] result543;
wire  [15:0] result544;
wire  [15:0] result545;
wire  [15:0] result546;
wire  [15:0] result547;
wire  [15:0] result548;
wire  [15:0] result549;
wire  [15:0] result550;
wire  [15:0] result551;
wire  [15:0] result552;
wire  [15:0] result553;
wire  [15:0] result554;
wire  [15:0] result555;
wire  [15:0] result556;
wire  [15:0] result557;
wire  [15:0] result558;
wire  [15:0] result559;
wire  [15:0] result560;
wire  [15:0] result561;
wire  [15:0] result562;
wire  [15:0] result563;
wire  [15:0] result564;
wire  [15:0] result565;
wire  [15:0] result566;
wire  [15:0] result567;
wire  [15:0] result568;
wire  [15:0] result569;
wire  [15:0] result570;
wire  [15:0] result571;
wire  [15:0] result572;
wire  [15:0] result573;
wire  [15:0] result574;
wire  [15:0] result575;
wire  [15:0] result576;
wire  [15:0] result577;
wire  [15:0] result578;
wire  [15:0] result579;
wire  [15:0] result580;
wire  [15:0] result581;
wire  [15:0] result582;
wire  [15:0] result583;
wire  [15:0] result584;
wire  [15:0] result585;
wire  [15:0] result586;
wire  [15:0] result587;
wire  [15:0] result588;
wire  [15:0] result589;
wire  [15:0] result590;
wire  [15:0] result591;
wire  [15:0] result592;
wire  [15:0] result593;
wire  [15:0] result594;
wire  [15:0] result595;
wire  [15:0] result596;
wire  [15:0] result597;
wire  [15:0] result598;
wire  [15:0] result599;
wire  [15:0] result600;
wire  [15:0] result601;
wire  [15:0] result602;
wire  [15:0] result603;
wire  [15:0] result604;
wire  [15:0] result605;
wire  [15:0] result606;
wire  [15:0] result607;
wire  [15:0] result608;
wire  [15:0] result609;
wire  [15:0] result610;
wire  [15:0] result611;
wire  [15:0] result612;
wire  [15:0] result613;
wire  [15:0] result614;
wire  [15:0] result615;
wire  [15:0] result616;
wire  [15:0] result617;
wire  [15:0] result618;
wire  [15:0] result619;
wire  [15:0] result620;
wire  [15:0] result621;
wire  [15:0] result622;
wire  [15:0] result623;
wire  [15:0] result624;
wire  [15:0] result625;
wire  [15:0] result626;
wire  [15:0] result627;
wire  [15:0] result628;
wire  [15:0] result629;
wire  [15:0] result630;
wire  [15:0] result631;
wire  [15:0] result632;
wire  [15:0] result633;
wire  [15:0] result634;
wire  [15:0] result635;
wire  [15:0] result636;
wire  [15:0] result637;
wire  [15:0] result638;
wire  [15:0] result639;
wire  [15:0] result640;
wire  [15:0] result641;
wire  [15:0] result642;
wire  [15:0] result643;
wire  [15:0] result644;
wire  [15:0] result645;
wire  [15:0] result646;
wire  [15:0] result647;
wire  [15:0] result648;
wire  [15:0] result649;
wire  [15:0] result650;
wire  [15:0] result651;
wire  [15:0] result652;
wire  [15:0] result653;
wire  [15:0] result654;
wire  [15:0] result655;
wire  [15:0] result656;
wire  [15:0] result657;
wire  [15:0] result658;
wire  [15:0] result659;
wire  [15:0] result660;
wire  [15:0] result661;
wire  [15:0] result662;
wire  [15:0] result663;
wire  [15:0] result664;
wire  [15:0] result665;
wire  [15:0] result666;
wire  [15:0] result667;
wire  [15:0] result668;
wire  [15:0] result669;
wire  [15:0] result670;
wire  [15:0] result671;
wire  [15:0] result672;
wire  [15:0] result673;
wire  [15:0] result674;
wire  [15:0] result675;
wire  [15:0] result676;
wire  [15:0] result677;
wire  [15:0] result678;
wire  [15:0] result679;
wire  [15:0] result680;
wire  [15:0] result681;
wire  [15:0] result682;
wire  [15:0] result683;
wire  [15:0] result684;
wire  [15:0] result685;
wire  [15:0] result686;
wire  [15:0] result687;
wire  [15:0] result688;
wire  [15:0] result689;
wire  [15:0] result690;
wire  [15:0] result691;
wire  [15:0] result692;
wire  [15:0] result693;
wire  [15:0] result694;
wire  [15:0] result695;
wire  [15:0] result696;
wire  [15:0] result697;
wire  [15:0] result698;
wire  [15:0] result699;
wire  [15:0] result700;
wire  [15:0] result701;
wire  [15:0] result702;
wire  [15:0] result703;
wire  [15:0] result704;
wire  [15:0] result705;
wire  [15:0] result706;
wire  [15:0] result707;
wire  [15:0] result708;
wire  [15:0] result709;
wire  [15:0] result710;
wire  [15:0] result711;
wire  [15:0] result712;
wire  [15:0] result713;
wire  [15:0] result714;
wire  [15:0] result715;
wire  [15:0] result716;
wire  [15:0] result717;
wire  [15:0] result718;
wire  [15:0] result719;
wire  [15:0] result720;
wire  [15:0] result721;
wire  [15:0] result722;
wire  [15:0] result723;
wire  [15:0] result724;
wire  [15:0] result725;
wire  [15:0] result726;
wire  [15:0] result727;
wire  [15:0] result728;
wire  [15:0] result729;
wire  [15:0] result730;
wire  [15:0] result731;
wire  [15:0] result732;
wire  [15:0] result733;
wire  [15:0] result734;
wire  [15:0] result735;
wire  [15:0] result736;
wire  [15:0] result737;
wire  [15:0] result738;
wire  [15:0] result739;
wire  [15:0] result740;
wire  [15:0] result741;
wire  [15:0] result742;
wire  [15:0] result743;
wire  [15:0] result744;
wire  [15:0] result745;
wire  [15:0] result746;
wire  [15:0] result747;
wire  [15:0] result748;
wire  [15:0] result749;
wire  [15:0] result750;
wire  [15:0] result751;
wire  [15:0] result752;
wire  [15:0] result753;
wire  [15:0] result754;
wire  [15:0] result755;
wire  [15:0] result756;
wire  [15:0] result757;
wire  [15:0] result758;
wire  [15:0] result759;
wire  [15:0] result760;
wire  [15:0] result761;
wire  [15:0] result762;
wire  [15:0] result763;
wire  [15:0] result764;
wire  [15:0] result765;
wire  [15:0] result766;
wire  [15:0] result767;
wire  [15:0] result768;
wire  [15:0] result769;
wire  [15:0] result770;
wire  [15:0] result771;
wire  [15:0] result772;
wire  [15:0] result773;
wire  [15:0] result774;
wire  [15:0] result775;
wire  [15:0] result776;
wire  [15:0] result777;
wire  [15:0] result778;
wire  [15:0] result779;
wire  [15:0] result780;
wire  [15:0] result781;
wire  [15:0] result782;
wire  [15:0] result783;
wire  [15:0] result784;
wire  [15:0] result785;
wire  [15:0] result786;
wire  [15:0] result787;
wire  [15:0] result788;
wire  [15:0] result789;
wire  [15:0] result790;
wire  [15:0] result791;
wire  [15:0] result792;
wire  [15:0] result793;
wire  [15:0] result794;
wire  [15:0] result795;
wire  [15:0] result796;
wire  [15:0] result797;
wire  [15:0] result798;
wire  [15:0] result799;
wire  [15:0] result800;
wire  [15:0] result801;
wire  [15:0] result802;
wire  [15:0] result803;
wire  [15:0] result804;
wire  [15:0] result805;
wire  [15:0] result806;
wire  [15:0] result807;
wire  [15:0] result808;
wire  [15:0] result809;
wire  [15:0] result810;
wire  [15:0] result811;
wire  [15:0] result812;
wire  [15:0] result813;
wire  [15:0] result814;
wire  [15:0] result815;
wire  [15:0] result816;
wire  [15:0] result817;
wire  [15:0] result818;
wire  [15:0] result819;
wire  [15:0] result820;
wire  [15:0] result821;
wire  [15:0] result822;
wire  [15:0] result823;
wire  [15:0] result824;
wire  [15:0] result825;
wire  [15:0] result826;
wire  [15:0] result827;
wire  [15:0] result828;
wire  [15:0] result829;
wire  [15:0] result830;
wire  [15:0] result831;
wire  [15:0] result832;
wire  [15:0] result833;
wire  [15:0] result834;
wire  [15:0] result835;
wire  [15:0] result836;
wire  [15:0] result837;
wire  [15:0] result838;
wire  [15:0] result839;
wire  [15:0] result840;
wire  [15:0] result841;
wire  [15:0] result842;
wire  [15:0] result843;
wire  [15:0] result844;
wire  [15:0] result845;
wire  [15:0] result846;
wire  [15:0] result847;
wire  [15:0] result848;
wire  [15:0] result849;
wire  [15:0] result850;
wire  [15:0] result851;
wire  [15:0] result852;
wire  [15:0] result853;
wire  [15:0] result854;
wire  [15:0] result855;
wire  [15:0] result856;
wire  [15:0] result857;
wire  [15:0] result858;
wire  [15:0] result859;
wire  [15:0] result860;
wire  [15:0] result861;
wire  [15:0] result862;
wire  [15:0] result863;
wire  [15:0] result864;
wire  [15:0] result865;
wire  [15:0] result866;
wire  [15:0] result867;
wire  [15:0] result868;
wire  [15:0] result869;
wire  [15:0] result870;
wire  [15:0] result871;
wire  [15:0] result872;
wire  [15:0] result873;
wire  [15:0] result874;
wire  [15:0] result875;
wire  [15:0] result876;
wire  [15:0] result877;
wire  [15:0] result878;
wire  [15:0] result879;
wire  [15:0] result880;
wire  [15:0] result881;
wire  [15:0] result882;
wire  [15:0] result883;
wire  [15:0] result884;
wire  [15:0] result885;
wire  [15:0] result886;
wire  [15:0] result887;
wire  [15:0] result888;
wire  [15:0] result889;
wire  [15:0] result890;
wire  [15:0] result891;
wire  [15:0] result892;
wire  [15:0] result893;
wire  [15:0] result894;
wire  [15:0] result895;
wire  [15:0] result896;
wire  [15:0] result897;
wire  [15:0] result898;
wire  [15:0] result899;
wire  [15:0] result900;
wire  [15:0] result901;
wire  [15:0] result902;
wire  [15:0] result903;
wire  [15:0] result904;
wire  [15:0] result905;
wire  [15:0] result906;
wire  [15:0] result907;
wire  [15:0] result908;
wire  [15:0] result909;
wire  [15:0] result910;
wire  [15:0] result911;
wire  [15:0] result912;
wire  [15:0] result913;
wire  [15:0] result914;
wire  [15:0] result915;
wire  [15:0] result916;
wire  [15:0] result917;
wire  [15:0] result918;
wire  [15:0] result919;
wire  [15:0] result920;
wire  [15:0] result921;
wire  [15:0] result922;
wire  [15:0] result923;
wire  [15:0] result924;
wire  [15:0] result925;
wire  [15:0] result926;
wire  [15:0] result927;
wire  [15:0] result928;
wire  [15:0] result929;
wire  [15:0] result930;
wire  [15:0] result931;
wire  [15:0] result932;
wire  [15:0] result933;
wire  [15:0] result934;
wire  [15:0] result935;
wire  [15:0] result936;
wire  [15:0] result937;
wire  [15:0] result938;
wire  [15:0] result939;
wire  [15:0] result940;
wire  [15:0] result941;
wire  [15:0] result942;
wire  [15:0] result943;
wire  [15:0] result944;
wire  [15:0] result945;
wire  [15:0] result946;
wire  [15:0] result947;
wire  [15:0] result948;
wire  [15:0] result949;
wire  [15:0] result950;
wire  [15:0] result951;
wire  [15:0] result952;
wire  [15:0] result953;
wire  [15:0] result954;
wire  [15:0] result955;
wire  [15:0] result956;
wire  [15:0] result957;
wire  [15:0] result958;
wire  [15:0] result959;
wire  [15:0] result960;
wire  [15:0] result961;
wire  [15:0] result962;
wire  [15:0] result963;
wire  [15:0] result964;
wire  [15:0] result965;
wire  [15:0] result966;
wire  [15:0] result967;
wire  [15:0] result968;
wire  [15:0] result969;
wire  [15:0] result970;
wire  [15:0] result971;
wire  [15:0] result972;
wire  [15:0] result973;
wire  [15:0] result974;
wire  [15:0] result975;
wire  [15:0] result976;
wire  [15:0] result977;
wire  [15:0] result978;
wire  [15:0] result979;
wire  [15:0] result980;
wire  [15:0] result981;
wire  [15:0] result982;
wire  [15:0] result983;
wire  [15:0] result984;
wire  [15:0] result985;
wire  [15:0] result986;
wire  [15:0] result987;
wire  [15:0] result988;
wire  [15:0] result989;
wire  [15:0] result990;
wire  [15:0] result991;
wire  [15:0] result992;
wire  [15:0] result993;
wire  [15:0] result994;
wire  [15:0] result995;
wire  [15:0] result996;
wire  [15:0] result997;
wire  [15:0] result998;
wire  [15:0] result999;
wire  [15:0] result1000;
wire  [15:0] result1001;
wire  [15:0] result1002;
wire  [15:0] result1003;
wire  [15:0] result1004;
wire  [15:0] result1005;
wire  [15:0] result1006;
wire  [15:0] result1007;
wire  [15:0] result1008;
wire  [15:0] result1009;
wire  [15:0] result1010;
wire  [15:0] result1011;
wire  [15:0] result1012;
wire  [15:0] result1013;
wire  [15:0] result1014;
wire  [15:0] result1015;
wire  [15:0] result1016;
wire  [15:0] result1017;
wire  [15:0] result1018;
wire  [15:0] result1019;
wire  [15:0] result1020;
wire  [15:0] result1021;
wire  [15:0] result1022;
wire  [15:0] result1023;

PE P0 (inp_n0, inp_w0, clk, rst, out_s0, out_e0, result0);

PE P1(inp_n1, out_e1, clk, rst, out_s1, out_e1, result1);
PE P2(inp_n2, out_e2, clk, rst, out_s2, out_e2, result2);
PE P3(inp_n3, out_e3, clk, rst, out_s3, out_e3, result3);
PE P4(inp_n4, out_e4, clk, rst, out_s4, out_e4, result4);
PE P5(inp_n5, out_e5, clk, rst, out_s5, out_e5, result5);
PE P6(inp_n6, out_e6, clk, rst, out_s6, out_e6, result6);
PE P7(inp_n7, out_e7, clk, rst, out_s7, out_e7, result7);
PE P8(inp_n8, out_e8, clk, rst, out_s8, out_e8, result8);
PE P9(inp_n9, out_e9, clk, rst, out_s9, out_e9, result9);
PE P10(inp_n10, out_e10, clk, rst, out_s10, out_e10, result10);
PE P11(inp_n11, out_e11, clk, rst, out_s11, out_e11, result11);
PE P12(inp_n12, out_e12, clk, rst, out_s12, out_e12, result12);
PE P13(inp_n13, out_e13, clk, rst, out_s13, out_e13, result13);
PE P14(inp_n14, out_e14, clk, rst, out_s14, out_e14, result14);
PE P15(inp_n15, out_e15, clk, rst, out_s15, out_e15, result15);
PE P16(inp_n16, out_e16, clk, rst, out_s16, out_e16, result16);
PE P17(inp_n17, out_e17, clk, rst, out_s17, out_e17, result17);
PE P18(inp_n18, out_e18, clk, rst, out_s18, out_e18, result18);
PE P19(inp_n19, out_e19, clk, rst, out_s19, out_e19, result19);
PE P20(inp_n20, out_e20, clk, rst, out_s20, out_e20, result20);
PE P21(inp_n21, out_e21, clk, rst, out_s21, out_e21, result21);
PE P22(inp_n22, out_e22, clk, rst, out_s22, out_e22, result22);
PE P23(inp_n23, out_e23, clk, rst, out_s23, out_e23, result23);
PE P24(inp_n24, out_e24, clk, rst, out_s24, out_e24, result24);
PE P25(inp_n25, out_e25, clk, rst, out_s25, out_e25, result25);
PE P26(inp_n26, out_e26, clk, rst, out_s26, out_e26, result26);
PE P27(inp_n27, out_e27, clk, rst, out_s27, out_e27, result27);
PE P28(inp_n28, out_e28, clk, rst, out_s28, out_e28, result28);
PE P29(inp_n29, out_e29, clk, rst, out_s29, out_e29, result29);
PE P30(inp_n30, out_e30, clk, rst, out_s30, out_e30, result30);
PE P31(inp_n31, out_e31, clk, rst, out_s31, out_e31, result31);

PE P32(out_s0, inp_w32, clk, rst, out_s32, out_e32, result32);
PE P64(out_s32, inp_w64, clk, rst, out_s64, out_e64, result64);
PE P96(out_s64, inp_w96, clk, rst, out_s96, out_e96, result96);
PE P128(out_s96, inp_w128, clk, rst, out_s128, out_e128, result128);
PE P160(out_s128, inp_w160, clk, rst, out_s160, out_e160, result160);
PE P192(out_s160, inp_w192, clk, rst, out_s192, out_e192, result192);
PE P224(out_s192, inp_w224, clk, rst, out_s224, out_e224, result224);
PE P256(out_s224, inp_w256, clk, rst, out_s256, out_e256, result256);
PE P288(out_s256, inp_w288, clk, rst, out_s288, out_e288, result288);
PE P320(out_s288, inp_w320, clk, rst, out_s320, out_e320, result320);
PE P352(out_s320, inp_w352, clk, rst, out_s352, out_e352, result352);
PE P384(out_s352, inp_w384, clk, rst, out_s384, out_e384, result384);
PE P416(out_s384, inp_w416, clk, rst, out_s416, out_e416, result416);
PE P448(out_s416, inp_w448, clk, rst, out_s448, out_e448, result448);
PE P480(out_s448, inp_w480, clk, rst, out_s480, out_e480, result480);
PE P512(out_s480, inp_w512, clk, rst, out_s512, out_e512, result512);
PE P544(out_s512, inp_w544, clk, rst, out_s544, out_e544, result544);
PE P576(out_s544, inp_w576, clk, rst, out_s576, out_e576, result576);
PE P608(out_s576, inp_w608, clk, rst, out_s608, out_e608, result608);
PE P640(out_s608, inp_w640, clk, rst, out_s640, out_e640, result640);
PE P672(out_s640, inp_w672, clk, rst, out_s672, out_e672, result672);
PE P704(out_s672, inp_w704, clk, rst, out_s704, out_e704, result704);
PE P736(out_s704, inp_w736, clk, rst, out_s736, out_e736, result736);
PE P768(out_s736, inp_w768, clk, rst, out_s768, out_e768, result768);
PE P800(out_s768, inp_w800, clk, rst, out_s800, out_e800, result800);
PE P832(out_s800, inp_w832, clk, rst, out_s832, out_e832, result832);
PE P864(out_s832, inp_w864, clk, rst, out_s864, out_e864, result864);
PE P896(out_s864, inp_w896, clk, rst, out_s896, out_e896, result896);
PE P928(out_s896, inp_w928, clk, rst, out_s928, out_e928, result928);
PE P960(out_s928, inp_w960, clk, rst, out_s960, out_e960, result960);
PE P992(out_s960, inp_w992, clk, rst, out_s992, out_e992, result992);

PE P33(out_s1, out_e32, clk, rst, out_s33, out_e33, result33);
PE P34(out_s2, out_e33, clk, rst, out_s34, out_e34, result34);
PE P35(out_s3, out_e34, clk, rst, out_s35, out_e35, result35);
PE P36(out_s4, out_e35, clk, rst, out_s36, out_e36, result36);
PE P37(out_s5, out_e36, clk, rst, out_s37, out_e37, result37);
PE P38(out_s6, out_e37, clk, rst, out_s38, out_e38, result38);
PE P39(out_s7, out_e38, clk, rst, out_s39, out_e39, result39);
PE P40(out_s8, out_e39, clk, rst, out_s40, out_e40, result40);
PE P41(out_s9, out_e40, clk, rst, out_s41, out_e41, result41);
PE P42(out_s10, out_e41, clk, rst, out_s42, out_e42, result42);
PE P43(out_s11, out_e42, clk, rst, out_s43, out_e43, result43);
PE P44(out_s12, out_e43, clk, rst, out_s44, out_e44, result44);
PE P45(out_s13, out_e44, clk, rst, out_s45, out_e45, result45);
PE P46(out_s14, out_e45, clk, rst, out_s46, out_e46, result46);
PE P47(out_s15, out_e46, clk, rst, out_s47, out_e47, result47);
PE P48(out_s16, out_e47, clk, rst, out_s48, out_e48, result48);
PE P49(out_s17, out_e48, clk, rst, out_s49, out_e49, result49);
PE P50(out_s18, out_e49, clk, rst, out_s50, out_e50, result50);
PE P51(out_s19, out_e50, clk, rst, out_s51, out_e51, result51);
PE P52(out_s20, out_e51, clk, rst, out_s52, out_e52, result52);
PE P53(out_s21, out_e52, clk, rst, out_s53, out_e53, result53);
PE P54(out_s22, out_e53, clk, rst, out_s54, out_e54, result54);
PE P55(out_s23, out_e54, clk, rst, out_s55, out_e55, result55);
PE P56(out_s24, out_e55, clk, rst, out_s56, out_e56, result56);
PE P57(out_s25, out_e56, clk, rst, out_s57, out_e57, result57);
PE P58(out_s26, out_e57, clk, rst, out_s58, out_e58, result58);
PE P59(out_s27, out_e58, clk, rst, out_s59, out_e59, result59);
PE P60(out_s28, out_e59, clk, rst, out_s60, out_e60, result60);
PE P61(out_s29, out_e60, clk, rst, out_s61, out_e61, result61);
PE P62(out_s30, out_e61, clk, rst, out_s62, out_e62, result62);
PE P63(out_s31, out_e62, clk, rst, out_s63, out_e63, result63);

PE P65(out_s33, out_e64, clk, rst, out_s65, out_e65, result65);
PE P66(out_s34, out_e65, clk, rst, out_s66, out_e66, result66);
PE P67(out_s35, out_e66, clk, rst, out_s67, out_e67, result67);
PE P68(out_s36, out_e67, clk, rst, out_s68, out_e68, result68);
PE P69(out_s37, out_e68, clk, rst, out_s69, out_e69, result69);
PE P70(out_s38, out_e69, clk, rst, out_s70, out_e70, result70);
PE P71(out_s39, out_e70, clk, rst, out_s71, out_e71, result71);
PE P72(out_s40, out_e71, clk, rst, out_s72, out_e72, result72);
PE P73(out_s41, out_e72, clk, rst, out_s73, out_e73, result73);
PE P74(out_s42, out_e73, clk, rst, out_s74, out_e74, result74);
PE P75(out_s43, out_e74, clk, rst, out_s75, out_e75, result75);
PE P76(out_s44, out_e75, clk, rst, out_s76, out_e76, result76);
PE P77(out_s45, out_e76, clk, rst, out_s77, out_e77, result77);
PE P78(out_s46, out_e77, clk, rst, out_s78, out_e78, result78);
PE P79(out_s47, out_e78, clk, rst, out_s79, out_e79, result79);
PE P80(out_s48, out_e79, clk, rst, out_s80, out_e80, result80);
PE P81(out_s49, out_e80, clk, rst, out_s81, out_e81, result81);
PE P82(out_s50, out_e81, clk, rst, out_s82, out_e82, result82);
PE P83(out_s51, out_e82, clk, rst, out_s83, out_e83, result83);
PE P84(out_s52, out_e83, clk, rst, out_s84, out_e84, result84);
PE P85(out_s53, out_e84, clk, rst, out_s85, out_e85, result85);
PE P86(out_s54, out_e85, clk, rst, out_s86, out_e86, result86);
PE P87(out_s55, out_e86, clk, rst, out_s87, out_e87, result87);
PE P88(out_s56, out_e87, clk, rst, out_s88, out_e88, result88);
PE P89(out_s57, out_e88, clk, rst, out_s89, out_e89, result89);
PE P90(out_s58, out_e89, clk, rst, out_s90, out_e90, result90);
PE P91(out_s59, out_e90, clk, rst, out_s91, out_e91, result91);
PE P92(out_s60, out_e91, clk, rst, out_s92, out_e92, result92);
PE P93(out_s61, out_e92, clk, rst, out_s93, out_e93, result93);
PE P94(out_s62, out_e93, clk, rst, out_s94, out_e94, result94);
PE P95(out_s63, out_e94, clk, rst, out_s95, out_e95, result95);

PE P97(out_s65, out_e96, clk, rst, out_s97, out_e97, result97);
PE P98(out_s66, out_e97, clk, rst, out_s98, out_e98, result98);
PE P99(out_s67, out_e98, clk, rst, out_s99, out_e99, result99);
PE P100(out_s68, out_e99, clk, rst, out_s100, out_e100, result100);
PE P101(out_s69, out_e100, clk, rst, out_s101, out_e101, result101);
PE P102(out_s70, out_e101, clk, rst, out_s102, out_e102, result102);
PE P103(out_s71, out_e102, clk, rst, out_s103, out_e103, result103);
PE P104(out_s72, out_e103, clk, rst, out_s104, out_e104, result104);
PE P105(out_s73, out_e104, clk, rst, out_s105, out_e105, result105);
PE P106(out_s74, out_e105, clk, rst, out_s106, out_e106, result106);
PE P107(out_s75, out_e106, clk, rst, out_s107, out_e107, result107);
PE P108(out_s76, out_e107, clk, rst, out_s108, out_e108, result108);
PE P109(out_s77, out_e108, clk, rst, out_s109, out_e109, result109);
PE P110(out_s78, out_e109, clk, rst, out_s110, out_e110, result110);
PE P111(out_s79, out_e110, clk, rst, out_s111, out_e111, result111);
PE P112(out_s80, out_e111, clk, rst, out_s112, out_e112, result112);
PE P113(out_s81, out_e112, clk, rst, out_s113, out_e113, result113);
PE P114(out_s82, out_e113, clk, rst, out_s114, out_e114, result114);
PE P115(out_s83, out_e114, clk, rst, out_s115, out_e115, result115);
PE P116(out_s84, out_e115, clk, rst, out_s116, out_e116, result116);
PE P117(out_s85, out_e116, clk, rst, out_s117, out_e117, result117);
PE P118(out_s86, out_e117, clk, rst, out_s118, out_e118, result118);
PE P119(out_s87, out_e118, clk, rst, out_s119, out_e119, result119);
PE P120(out_s88, out_e119, clk, rst, out_s120, out_e120, result120);
PE P121(out_s89, out_e120, clk, rst, out_s121, out_e121, result121);
PE P122(out_s90, out_e121, clk, rst, out_s122, out_e122, result122);
PE P123(out_s91, out_e122, clk, rst, out_s123, out_e123, result123);
PE P124(out_s92, out_e123, clk, rst, out_s124, out_e124, result124);
PE P125(out_s93, out_e124, clk, rst, out_s125, out_e125, result125);
PE P126(out_s94, out_e125, clk, rst, out_s126, out_e126, result126);
PE P127(out_s95, out_e126, clk, rst, out_s127, out_e127, result127);

PE P129(out_s97, out_e128, clk, rst, out_s129, out_e129, result129);
PE P130(out_s98, out_e129, clk, rst, out_s130, out_e130, result130);
PE P131(out_s99, out_e130, clk, rst, out_s131, out_e131, result131);
PE P132(out_s100, out_e131, clk, rst, out_s132, out_e132, result132);
PE P133(out_s101, out_e132, clk, rst, out_s133, out_e133, result133);
PE P134(out_s102, out_e133, clk, rst, out_s134, out_e134, result134);
PE P135(out_s103, out_e134, clk, rst, out_s135, out_e135, result135);
PE P136(out_s104, out_e135, clk, rst, out_s136, out_e136, result136);
PE P137(out_s105, out_e136, clk, rst, out_s137, out_e137, result137);
PE P138(out_s106, out_e137, clk, rst, out_s138, out_e138, result138);
PE P139(out_s107, out_e138, clk, rst, out_s139, out_e139, result139);
PE P140(out_s108, out_e139, clk, rst, out_s140, out_e140, result140);
PE P141(out_s109, out_e140, clk, rst, out_s141, out_e141, result141);
PE P142(out_s110, out_e141, clk, rst, out_s142, out_e142, result142);
PE P143(out_s111, out_e142, clk, rst, out_s143, out_e143, result143);
PE P144(out_s112, out_e143, clk, rst, out_s144, out_e144, result144);
PE P145(out_s113, out_e144, clk, rst, out_s145, out_e145, result145);
PE P146(out_s114, out_e145, clk, rst, out_s146, out_e146, result146);
PE P147(out_s115, out_e146, clk, rst, out_s147, out_e147, result147);
PE P148(out_s116, out_e147, clk, rst, out_s148, out_e148, result148);
PE P149(out_s117, out_e148, clk, rst, out_s149, out_e149, result149);
PE P150(out_s118, out_e149, clk, rst, out_s150, out_e150, result150);
PE P151(out_s119, out_e150, clk, rst, out_s151, out_e151, result151);
PE P152(out_s120, out_e151, clk, rst, out_s152, out_e152, result152);
PE P153(out_s121, out_e152, clk, rst, out_s153, out_e153, result153);
PE P154(out_s122, out_e153, clk, rst, out_s154, out_e154, result154);
PE P155(out_s123, out_e154, clk, rst, out_s155, out_e155, result155);
PE P156(out_s124, out_e155, clk, rst, out_s156, out_e156, result156);
PE P157(out_s125, out_e156, clk, rst, out_s157, out_e157, result157);
PE P158(out_s126, out_e157, clk, rst, out_s158, out_e158, result158);
PE P159(out_s127, out_e158, clk, rst, out_s159, out_e159, result159);

PE P161(out_s129, out_e160, clk, rst, out_s161, out_e161, result161);
PE P162(out_s130, out_e161, clk, rst, out_s162, out_e162, result162);
PE P163(out_s131, out_e162, clk, rst, out_s163, out_e163, result163);
PE P164(out_s132, out_e163, clk, rst, out_s164, out_e164, result164);
PE P165(out_s133, out_e164, clk, rst, out_s165, out_e165, result165);
PE P166(out_s134, out_e165, clk, rst, out_s166, out_e166, result166);
PE P167(out_s135, out_e166, clk, rst, out_s167, out_e167, result167);
PE P168(out_s136, out_e167, clk, rst, out_s168, out_e168, result168);
PE P169(out_s137, out_e168, clk, rst, out_s169, out_e169, result169);
PE P170(out_s138, out_e169, clk, rst, out_s170, out_e170, result170);
PE P171(out_s139, out_e170, clk, rst, out_s171, out_e171, result171);
PE P172(out_s140, out_e171, clk, rst, out_s172, out_e172, result172);
PE P173(out_s141, out_e172, clk, rst, out_s173, out_e173, result173);
PE P174(out_s142, out_e173, clk, rst, out_s174, out_e174, result174);
PE P175(out_s143, out_e174, clk, rst, out_s175, out_e175, result175);
PE P176(out_s144, out_e175, clk, rst, out_s176, out_e176, result176);
PE P177(out_s145, out_e176, clk, rst, out_s177, out_e177, result177);
PE P178(out_s146, out_e177, clk, rst, out_s178, out_e178, result178);
PE P179(out_s147, out_e178, clk, rst, out_s179, out_e179, result179);
PE P180(out_s148, out_e179, clk, rst, out_s180, out_e180, result180);
PE P181(out_s149, out_e180, clk, rst, out_s181, out_e181, result181);
PE P182(out_s150, out_e181, clk, rst, out_s182, out_e182, result182);
PE P183(out_s151, out_e182, clk, rst, out_s183, out_e183, result183);
PE P184(out_s152, out_e183, clk, rst, out_s184, out_e184, result184);
PE P185(out_s153, out_e184, clk, rst, out_s185, out_e185, result185);
PE P186(out_s154, out_e185, clk, rst, out_s186, out_e186, result186);
PE P187(out_s155, out_e186, clk, rst, out_s187, out_e187, result187);
PE P188(out_s156, out_e187, clk, rst, out_s188, out_e188, result188);
PE P189(out_s157, out_e188, clk, rst, out_s189, out_e189, result189);
PE P190(out_s158, out_e189, clk, rst, out_s190, out_e190, result190);
PE P191(out_s159, out_e190, clk, rst, out_s191, out_e191, result191);

PE P193(out_s161, out_e192, clk, rst, out_s193, out_e193, result193);
PE P194(out_s162, out_e193, clk, rst, out_s194, out_e194, result194);
PE P195(out_s163, out_e194, clk, rst, out_s195, out_e195, result195);
PE P196(out_s164, out_e195, clk, rst, out_s196, out_e196, result196);
PE P197(out_s165, out_e196, clk, rst, out_s197, out_e197, result197);
PE P198(out_s166, out_e197, clk, rst, out_s198, out_e198, result198);
PE P199(out_s167, out_e198, clk, rst, out_s199, out_e199, result199);
PE P200(out_s168, out_e199, clk, rst, out_s200, out_e200, result200);
PE P201(out_s169, out_e200, clk, rst, out_s201, out_e201, result201);
PE P202(out_s170, out_e201, clk, rst, out_s202, out_e202, result202);
PE P203(out_s171, out_e202, clk, rst, out_s203, out_e203, result203);
PE P204(out_s172, out_e203, clk, rst, out_s204, out_e204, result204);
PE P205(out_s173, out_e204, clk, rst, out_s205, out_e205, result205);
PE P206(out_s174, out_e205, clk, rst, out_s206, out_e206, result206);
PE P207(out_s175, out_e206, clk, rst, out_s207, out_e207, result207);
PE P208(out_s176, out_e207, clk, rst, out_s208, out_e208, result208);
PE P209(out_s177, out_e208, clk, rst, out_s209, out_e209, result209);
PE P210(out_s178, out_e209, clk, rst, out_s210, out_e210, result210);
PE P211(out_s179, out_e210, clk, rst, out_s211, out_e211, result211);
PE P212(out_s180, out_e211, clk, rst, out_s212, out_e212, result212);
PE P213(out_s181, out_e212, clk, rst, out_s213, out_e213, result213);
PE P214(out_s182, out_e213, clk, rst, out_s214, out_e214, result214);
PE P215(out_s183, out_e214, clk, rst, out_s215, out_e215, result215);
PE P216(out_s184, out_e215, clk, rst, out_s216, out_e216, result216);
PE P217(out_s185, out_e216, clk, rst, out_s217, out_e217, result217);
PE P218(out_s186, out_e217, clk, rst, out_s218, out_e218, result218);
PE P219(out_s187, out_e218, clk, rst, out_s219, out_e219, result219);
PE P220(out_s188, out_e219, clk, rst, out_s220, out_e220, result220);
PE P221(out_s189, out_e220, clk, rst, out_s221, out_e221, result221);
PE P222(out_s190, out_e221, clk, rst, out_s222, out_e222, result222);
PE P223(out_s191, out_e222, clk, rst, out_s223, out_e223, result223);

PE P225(out_s193, out_e224, clk, rst, out_s225, out_e225, result225);
PE P226(out_s194, out_e225, clk, rst, out_s226, out_e226, result226);
PE P227(out_s195, out_e226, clk, rst, out_s227, out_e227, result227);
PE P228(out_s196, out_e227, clk, rst, out_s228, out_e228, result228);
PE P229(out_s197, out_e228, clk, rst, out_s229, out_e229, result229);
PE P230(out_s198, out_e229, clk, rst, out_s230, out_e230, result230);
PE P231(out_s199, out_e230, clk, rst, out_s231, out_e231, result231);
PE P232(out_s200, out_e231, clk, rst, out_s232, out_e232, result232);
PE P233(out_s201, out_e232, clk, rst, out_s233, out_e233, result233);
PE P234(out_s202, out_e233, clk, rst, out_s234, out_e234, result234);
PE P235(out_s203, out_e234, clk, rst, out_s235, out_e235, result235);
PE P236(out_s204, out_e235, clk, rst, out_s236, out_e236, result236);
PE P237(out_s205, out_e236, clk, rst, out_s237, out_e237, result237);
PE P238(out_s206, out_e237, clk, rst, out_s238, out_e238, result238);
PE P239(out_s207, out_e238, clk, rst, out_s239, out_e239, result239);
PE P240(out_s208, out_e239, clk, rst, out_s240, out_e240, result240);
PE P241(out_s209, out_e240, clk, rst, out_s241, out_e241, result241);
PE P242(out_s210, out_e241, clk, rst, out_s242, out_e242, result242);
PE P243(out_s211, out_e242, clk, rst, out_s243, out_e243, result243);
PE P244(out_s212, out_e243, clk, rst, out_s244, out_e244, result244);
PE P245(out_s213, out_e244, clk, rst, out_s245, out_e245, result245);
PE P246(out_s214, out_e245, clk, rst, out_s246, out_e246, result246);
PE P247(out_s215, out_e246, clk, rst, out_s247, out_e247, result247);
PE P248(out_s216, out_e247, clk, rst, out_s248, out_e248, result248);
PE P249(out_s217, out_e248, clk, rst, out_s249, out_e249, result249);
PE P250(out_s218, out_e249, clk, rst, out_s250, out_e250, result250);
PE P251(out_s219, out_e250, clk, rst, out_s251, out_e251, result251);
PE P252(out_s220, out_e251, clk, rst, out_s252, out_e252, result252);
PE P253(out_s221, out_e252, clk, rst, out_s253, out_e253, result253);
PE P254(out_s222, out_e253, clk, rst, out_s254, out_e254, result254);
PE P255(out_s223, out_e254, clk, rst, out_s255, out_e255, result255);

PE P257(out_s225, out_e256, clk, rst, out_s257, out_e257, result257);
PE P258(out_s226, out_e257, clk, rst, out_s258, out_e258, result258);
PE P259(out_s227, out_e258, clk, rst, out_s259, out_e259, result259);
PE P260(out_s228, out_e259, clk, rst, out_s260, out_e260, result260);
PE P261(out_s229, out_e260, clk, rst, out_s261, out_e261, result261);
PE P262(out_s230, out_e261, clk, rst, out_s262, out_e262, result262);
PE P263(out_s231, out_e262, clk, rst, out_s263, out_e263, result263);
PE P264(out_s232, out_e263, clk, rst, out_s264, out_e264, result264);
PE P265(out_s233, out_e264, clk, rst, out_s265, out_e265, result265);
PE P266(out_s234, out_e265, clk, rst, out_s266, out_e266, result266);
PE P267(out_s235, out_e266, clk, rst, out_s267, out_e267, result267);
PE P268(out_s236, out_e267, clk, rst, out_s268, out_e268, result268);
PE P269(out_s237, out_e268, clk, rst, out_s269, out_e269, result269);
PE P270(out_s238, out_e269, clk, rst, out_s270, out_e270, result270);
PE P271(out_s239, out_e270, clk, rst, out_s271, out_e271, result271);
PE P272(out_s240, out_e271, clk, rst, out_s272, out_e272, result272);
PE P273(out_s241, out_e272, clk, rst, out_s273, out_e273, result273);
PE P274(out_s242, out_e273, clk, rst, out_s274, out_e274, result274);
PE P275(out_s243, out_e274, clk, rst, out_s275, out_e275, result275);
PE P276(out_s244, out_e275, clk, rst, out_s276, out_e276, result276);
PE P277(out_s245, out_e276, clk, rst, out_s277, out_e277, result277);
PE P278(out_s246, out_e277, clk, rst, out_s278, out_e278, result278);
PE P279(out_s247, out_e278, clk, rst, out_s279, out_e279, result279);
PE P280(out_s248, out_e279, clk, rst, out_s280, out_e280, result280);
PE P281(out_s249, out_e280, clk, rst, out_s281, out_e281, result281);
PE P282(out_s250, out_e281, clk, rst, out_s282, out_e282, result282);
PE P283(out_s251, out_e282, clk, rst, out_s283, out_e283, result283);
PE P284(out_s252, out_e283, clk, rst, out_s284, out_e284, result284);
PE P285(out_s253, out_e284, clk, rst, out_s285, out_e285, result285);
PE P286(out_s254, out_e285, clk, rst, out_s286, out_e286, result286);
PE P287(out_s255, out_e286, clk, rst, out_s287, out_e287, result287);

PE P289(out_s257, out_e288, clk, rst, out_s289, out_e289, result289);
PE P290(out_s258, out_e289, clk, rst, out_s290, out_e290, result290);
PE P291(out_s259, out_e290, clk, rst, out_s291, out_e291, result291);
PE P292(out_s260, out_e291, clk, rst, out_s292, out_e292, result292);
PE P293(out_s261, out_e292, clk, rst, out_s293, out_e293, result293);
PE P294(out_s262, out_e293, clk, rst, out_s294, out_e294, result294);
PE P295(out_s263, out_e294, clk, rst, out_s295, out_e295, result295);
PE P296(out_s264, out_e295, clk, rst, out_s296, out_e296, result296);
PE P297(out_s265, out_e296, clk, rst, out_s297, out_e297, result297);
PE P298(out_s266, out_e297, clk, rst, out_s298, out_e298, result298);
PE P299(out_s267, out_e298, clk, rst, out_s299, out_e299, result299);
PE P300(out_s268, out_e299, clk, rst, out_s300, out_e300, result300);
PE P301(out_s269, out_e300, clk, rst, out_s301, out_e301, result301);
PE P302(out_s270, out_e301, clk, rst, out_s302, out_e302, result302);
PE P303(out_s271, out_e302, clk, rst, out_s303, out_e303, result303);
PE P304(out_s272, out_e303, clk, rst, out_s304, out_e304, result304);
PE P305(out_s273, out_e304, clk, rst, out_s305, out_e305, result305);
PE P306(out_s274, out_e305, clk, rst, out_s306, out_e306, result306);
PE P307(out_s275, out_e306, clk, rst, out_s307, out_e307, result307);
PE P308(out_s276, out_e307, clk, rst, out_s308, out_e308, result308);
PE P309(out_s277, out_e308, clk, rst, out_s309, out_e309, result309);
PE P310(out_s278, out_e309, clk, rst, out_s310, out_e310, result310);
PE P311(out_s279, out_e310, clk, rst, out_s311, out_e311, result311);
PE P312(out_s280, out_e311, clk, rst, out_s312, out_e312, result312);
PE P313(out_s281, out_e312, clk, rst, out_s313, out_e313, result313);
PE P314(out_s282, out_e313, clk, rst, out_s314, out_e314, result314);
PE P315(out_s283, out_e314, clk, rst, out_s315, out_e315, result315);
PE P316(out_s284, out_e315, clk, rst, out_s316, out_e316, result316);
PE P317(out_s285, out_e316, clk, rst, out_s317, out_e317, result317);
PE P318(out_s286, out_e317, clk, rst, out_s318, out_e318, result318);
PE P319(out_s287, out_e318, clk, rst, out_s319, out_e319, result319);

PE P321(out_s289, out_e320, clk, rst, out_s321, out_e321, result321);
PE P322(out_s290, out_e321, clk, rst, out_s322, out_e322, result322);
PE P323(out_s291, out_e322, clk, rst, out_s323, out_e323, result323);
PE P324(out_s292, out_e323, clk, rst, out_s324, out_e324, result324);
PE P325(out_s293, out_e324, clk, rst, out_s325, out_e325, result325);
PE P326(out_s294, out_e325, clk, rst, out_s326, out_e326, result326);
PE P327(out_s295, out_e326, clk, rst, out_s327, out_e327, result327);
PE P328(out_s296, out_e327, clk, rst, out_s328, out_e328, result328);
PE P329(out_s297, out_e328, clk, rst, out_s329, out_e329, result329);
PE P330(out_s298, out_e329, clk, rst, out_s330, out_e330, result330);
PE P331(out_s299, out_e330, clk, rst, out_s331, out_e331, result331);
PE P332(out_s300, out_e331, clk, rst, out_s332, out_e332, result332);
PE P333(out_s301, out_e332, clk, rst, out_s333, out_e333, result333);
PE P334(out_s302, out_e333, clk, rst, out_s334, out_e334, result334);
PE P335(out_s303, out_e334, clk, rst, out_s335, out_e335, result335);
PE P336(out_s304, out_e335, clk, rst, out_s336, out_e336, result336);
PE P337(out_s305, out_e336, clk, rst, out_s337, out_e337, result337);
PE P338(out_s306, out_e337, clk, rst, out_s338, out_e338, result338);
PE P339(out_s307, out_e338, clk, rst, out_s339, out_e339, result339);
PE P340(out_s308, out_e339, clk, rst, out_s340, out_e340, result340);
PE P341(out_s309, out_e340, clk, rst, out_s341, out_e341, result341);
PE P342(out_s310, out_e341, clk, rst, out_s342, out_e342, result342);
PE P343(out_s311, out_e342, clk, rst, out_s343, out_e343, result343);
PE P344(out_s312, out_e343, clk, rst, out_s344, out_e344, result344);
PE P345(out_s313, out_e344, clk, rst, out_s345, out_e345, result345);
PE P346(out_s314, out_e345, clk, rst, out_s346, out_e346, result346);
PE P347(out_s315, out_e346, clk, rst, out_s347, out_e347, result347);
PE P348(out_s316, out_e347, clk, rst, out_s348, out_e348, result348);
PE P349(out_s317, out_e348, clk, rst, out_s349, out_e349, result349);
PE P350(out_s318, out_e349, clk, rst, out_s350, out_e350, result350);
PE P351(out_s319, out_e350, clk, rst, out_s351, out_e351, result351);

PE P353(out_s321, out_e352, clk, rst, out_s353, out_e353, result353);
PE P354(out_s322, out_e353, clk, rst, out_s354, out_e354, result354);
PE P355(out_s323, out_e354, clk, rst, out_s355, out_e355, result355);
PE P356(out_s324, out_e355, clk, rst, out_s356, out_e356, result356);
PE P357(out_s325, out_e356, clk, rst, out_s357, out_e357, result357);
PE P358(out_s326, out_e357, clk, rst, out_s358, out_e358, result358);
PE P359(out_s327, out_e358, clk, rst, out_s359, out_e359, result359);
PE P360(out_s328, out_e359, clk, rst, out_s360, out_e360, result360);
PE P361(out_s329, out_e360, clk, rst, out_s361, out_e361, result361);
PE P362(out_s330, out_e361, clk, rst, out_s362, out_e362, result362);
PE P363(out_s331, out_e362, clk, rst, out_s363, out_e363, result363);
PE P364(out_s332, out_e363, clk, rst, out_s364, out_e364, result364);
PE P365(out_s333, out_e364, clk, rst, out_s365, out_e365, result365);
PE P366(out_s334, out_e365, clk, rst, out_s366, out_e366, result366);
PE P367(out_s335, out_e366, clk, rst, out_s367, out_e367, result367);
PE P368(out_s336, out_e367, clk, rst, out_s368, out_e368, result368);
PE P369(out_s337, out_e368, clk, rst, out_s369, out_e369, result369);
PE P370(out_s338, out_e369, clk, rst, out_s370, out_e370, result370);
PE P371(out_s339, out_e370, clk, rst, out_s371, out_e371, result371);
PE P372(out_s340, out_e371, clk, rst, out_s372, out_e372, result372);
PE P373(out_s341, out_e372, clk, rst, out_s373, out_e373, result373);
PE P374(out_s342, out_e373, clk, rst, out_s374, out_e374, result374);
PE P375(out_s343, out_e374, clk, rst, out_s375, out_e375, result375);
PE P376(out_s344, out_e375, clk, rst, out_s376, out_e376, result376);
PE P377(out_s345, out_e376, clk, rst, out_s377, out_e377, result377);
PE P378(out_s346, out_e377, clk, rst, out_s378, out_e378, result378);
PE P379(out_s347, out_e378, clk, rst, out_s379, out_e379, result379);
PE P380(out_s348, out_e379, clk, rst, out_s380, out_e380, result380);
PE P381(out_s349, out_e380, clk, rst, out_s381, out_e381, result381);
PE P382(out_s350, out_e381, clk, rst, out_s382, out_e382, result382);
PE P383(out_s351, out_e382, clk, rst, out_s383, out_e383, result383);

PE P385(out_s353, out_e384, clk, rst, out_s385, out_e385, result385);
PE P386(out_s354, out_e385, clk, rst, out_s386, out_e386, result386);
PE P387(out_s355, out_e386, clk, rst, out_s387, out_e387, result387);
PE P388(out_s356, out_e387, clk, rst, out_s388, out_e388, result388);
PE P389(out_s357, out_e388, clk, rst, out_s389, out_e389, result389);
PE P390(out_s358, out_e389, clk, rst, out_s390, out_e390, result390);
PE P391(out_s359, out_e390, clk, rst, out_s391, out_e391, result391);
PE P392(out_s360, out_e391, clk, rst, out_s392, out_e392, result392);
PE P393(out_s361, out_e392, clk, rst, out_s393, out_e393, result393);
PE P394(out_s362, out_e393, clk, rst, out_s394, out_e394, result394);
PE P395(out_s363, out_e394, clk, rst, out_s395, out_e395, result395);
PE P396(out_s364, out_e395, clk, rst, out_s396, out_e396, result396);
PE P397(out_s365, out_e396, clk, rst, out_s397, out_e397, result397);
PE P398(out_s366, out_e397, clk, rst, out_s398, out_e398, result398);
PE P399(out_s367, out_e398, clk, rst, out_s399, out_e399, result399);
PE P400(out_s368, out_e399, clk, rst, out_s400, out_e400, result400);
PE P401(out_s369, out_e400, clk, rst, out_s401, out_e401, result401);
PE P402(out_s370, out_e401, clk, rst, out_s402, out_e402, result402);
PE P403(out_s371, out_e402, clk, rst, out_s403, out_e403, result403);
PE P404(out_s372, out_e403, clk, rst, out_s404, out_e404, result404);
PE P405(out_s373, out_e404, clk, rst, out_s405, out_e405, result405);
PE P406(out_s374, out_e405, clk, rst, out_s406, out_e406, result406);
PE P407(out_s375, out_e406, clk, rst, out_s407, out_e407, result407);
PE P408(out_s376, out_e407, clk, rst, out_s408, out_e408, result408);
PE P409(out_s377, out_e408, clk, rst, out_s409, out_e409, result409);
PE P410(out_s378, out_e409, clk, rst, out_s410, out_e410, result410);
PE P411(out_s379, out_e410, clk, rst, out_s411, out_e411, result411);
PE P412(out_s380, out_e411, clk, rst, out_s412, out_e412, result412);
PE P413(out_s381, out_e412, clk, rst, out_s413, out_e413, result413);
PE P414(out_s382, out_e413, clk, rst, out_s414, out_e414, result414);
PE P415(out_s383, out_e414, clk, rst, out_s415, out_e415, result415);

PE P417(out_s385, out_e416, clk, rst, out_s417, out_e417, result417);
PE P418(out_s386, out_e417, clk, rst, out_s418, out_e418, result418);
PE P419(out_s387, out_e418, clk, rst, out_s419, out_e419, result419);
PE P420(out_s388, out_e419, clk, rst, out_s420, out_e420, result420);
PE P421(out_s389, out_e420, clk, rst, out_s421, out_e421, result421);
PE P422(out_s390, out_e421, clk, rst, out_s422, out_e422, result422);
PE P423(out_s391, out_e422, clk, rst, out_s423, out_e423, result423);
PE P424(out_s392, out_e423, clk, rst, out_s424, out_e424, result424);
PE P425(out_s393, out_e424, clk, rst, out_s425, out_e425, result425);
PE P426(out_s394, out_e425, clk, rst, out_s426, out_e426, result426);
PE P427(out_s395, out_e426, clk, rst, out_s427, out_e427, result427);
PE P428(out_s396, out_e427, clk, rst, out_s428, out_e428, result428);
PE P429(out_s397, out_e428, clk, rst, out_s429, out_e429, result429);
PE P430(out_s398, out_e429, clk, rst, out_s430, out_e430, result430);
PE P431(out_s399, out_e430, clk, rst, out_s431, out_e431, result431);
PE P432(out_s400, out_e431, clk, rst, out_s432, out_e432, result432);
PE P433(out_s401, out_e432, clk, rst, out_s433, out_e433, result433);
PE P434(out_s402, out_e433, clk, rst, out_s434, out_e434, result434);
PE P435(out_s403, out_e434, clk, rst, out_s435, out_e435, result435);
PE P436(out_s404, out_e435, clk, rst, out_s436, out_e436, result436);
PE P437(out_s405, out_e436, clk, rst, out_s437, out_e437, result437);
PE P438(out_s406, out_e437, clk, rst, out_s438, out_e438, result438);
PE P439(out_s407, out_e438, clk, rst, out_s439, out_e439, result439);
PE P440(out_s408, out_e439, clk, rst, out_s440, out_e440, result440);
PE P441(out_s409, out_e440, clk, rst, out_s441, out_e441, result441);
PE P442(out_s410, out_e441, clk, rst, out_s442, out_e442, result442);
PE P443(out_s411, out_e442, clk, rst, out_s443, out_e443, result443);
PE P444(out_s412, out_e443, clk, rst, out_s444, out_e444, result444);
PE P445(out_s413, out_e444, clk, rst, out_s445, out_e445, result445);
PE P446(out_s414, out_e445, clk, rst, out_s446, out_e446, result446);
PE P447(out_s415, out_e446, clk, rst, out_s447, out_e447, result447);

PE P449(out_s417, out_e448, clk, rst, out_s449, out_e449, result449);
PE P450(out_s418, out_e449, clk, rst, out_s450, out_e450, result450);
PE P451(out_s419, out_e450, clk, rst, out_s451, out_e451, result451);
PE P452(out_s420, out_e451, clk, rst, out_s452, out_e452, result452);
PE P453(out_s421, out_e452, clk, rst, out_s453, out_e453, result453);
PE P454(out_s422, out_e453, clk, rst, out_s454, out_e454, result454);
PE P455(out_s423, out_e454, clk, rst, out_s455, out_e455, result455);
PE P456(out_s424, out_e455, clk, rst, out_s456, out_e456, result456);
PE P457(out_s425, out_e456, clk, rst, out_s457, out_e457, result457);
PE P458(out_s426, out_e457, clk, rst, out_s458, out_e458, result458);
PE P459(out_s427, out_e458, clk, rst, out_s459, out_e459, result459);
PE P460(out_s428, out_e459, clk, rst, out_s460, out_e460, result460);
PE P461(out_s429, out_e460, clk, rst, out_s461, out_e461, result461);
PE P462(out_s430, out_e461, clk, rst, out_s462, out_e462, result462);
PE P463(out_s431, out_e462, clk, rst, out_s463, out_e463, result463);
PE P464(out_s432, out_e463, clk, rst, out_s464, out_e464, result464);
PE P465(out_s433, out_e464, clk, rst, out_s465, out_e465, result465);
PE P466(out_s434, out_e465, clk, rst, out_s466, out_e466, result466);
PE P467(out_s435, out_e466, clk, rst, out_s467, out_e467, result467);
PE P468(out_s436, out_e467, clk, rst, out_s468, out_e468, result468);
PE P469(out_s437, out_e468, clk, rst, out_s469, out_e469, result469);
PE P470(out_s438, out_e469, clk, rst, out_s470, out_e470, result470);
PE P471(out_s439, out_e470, clk, rst, out_s471, out_e471, result471);
PE P472(out_s440, out_e471, clk, rst, out_s472, out_e472, result472);
PE P473(out_s441, out_e472, clk, rst, out_s473, out_e473, result473);
PE P474(out_s442, out_e473, clk, rst, out_s474, out_e474, result474);
PE P475(out_s443, out_e474, clk, rst, out_s475, out_e475, result475);
PE P476(out_s444, out_e475, clk, rst, out_s476, out_e476, result476);
PE P477(out_s445, out_e476, clk, rst, out_s477, out_e477, result477);
PE P478(out_s446, out_e477, clk, rst, out_s478, out_e478, result478);
PE P479(out_s447, out_e478, clk, rst, out_s479, out_e479, result479);

PE P481(out_s449, out_e480, clk, rst, out_s481, out_e481, result481);
PE P482(out_s450, out_e481, clk, rst, out_s482, out_e482, result482);
PE P483(out_s451, out_e482, clk, rst, out_s483, out_e483, result483);
PE P484(out_s452, out_e483, clk, rst, out_s484, out_e484, result484);
PE P485(out_s453, out_e484, clk, rst, out_s485, out_e485, result485);
PE P486(out_s454, out_e485, clk, rst, out_s486, out_e486, result486);
PE P487(out_s455, out_e486, clk, rst, out_s487, out_e487, result487);
PE P488(out_s456, out_e487, clk, rst, out_s488, out_e488, result488);
PE P489(out_s457, out_e488, clk, rst, out_s489, out_e489, result489);
PE P490(out_s458, out_e489, clk, rst, out_s490, out_e490, result490);
PE P491(out_s459, out_e490, clk, rst, out_s491, out_e491, result491);
PE P492(out_s460, out_e491, clk, rst, out_s492, out_e492, result492);
PE P493(out_s461, out_e492, clk, rst, out_s493, out_e493, result493);
PE P494(out_s462, out_e493, clk, rst, out_s494, out_e494, result494);
PE P495(out_s463, out_e494, clk, rst, out_s495, out_e495, result495);
PE P496(out_s464, out_e495, clk, rst, out_s496, out_e496, result496);
PE P497(out_s465, out_e496, clk, rst, out_s497, out_e497, result497);
PE P498(out_s466, out_e497, clk, rst, out_s498, out_e498, result498);
PE P499(out_s467, out_e498, clk, rst, out_s499, out_e499, result499);
PE P500(out_s468, out_e499, clk, rst, out_s500, out_e500, result500);
PE P501(out_s469, out_e500, clk, rst, out_s501, out_e501, result501);
PE P502(out_s470, out_e501, clk, rst, out_s502, out_e502, result502);
PE P503(out_s471, out_e502, clk, rst, out_s503, out_e503, result503);
PE P504(out_s472, out_e503, clk, rst, out_s504, out_e504, result504);
PE P505(out_s473, out_e504, clk, rst, out_s505, out_e505, result505);
PE P506(out_s474, out_e505, clk, rst, out_s506, out_e506, result506);
PE P507(out_s475, out_e506, clk, rst, out_s507, out_e507, result507);
PE P508(out_s476, out_e507, clk, rst, out_s508, out_e508, result508);
PE P509(out_s477, out_e508, clk, rst, out_s509, out_e509, result509);
PE P510(out_s478, out_e509, clk, rst, out_s510, out_e510, result510);
PE P511(out_s479, out_e510, clk, rst, out_s511, out_e511, result511);

PE P513(out_s481, out_e512, clk, rst, out_s513, out_e513, result513);
PE P514(out_s482, out_e513, clk, rst, out_s514, out_e514, result514);
PE P515(out_s483, out_e514, clk, rst, out_s515, out_e515, result515);
PE P516(out_s484, out_e515, clk, rst, out_s516, out_e516, result516);
PE P517(out_s485, out_e516, clk, rst, out_s517, out_e517, result517);
PE P518(out_s486, out_e517, clk, rst, out_s518, out_e518, result518);
PE P519(out_s487, out_e518, clk, rst, out_s519, out_e519, result519);
PE P520(out_s488, out_e519, clk, rst, out_s520, out_e520, result520);
PE P521(out_s489, out_e520, clk, rst, out_s521, out_e521, result521);
PE P522(out_s490, out_e521, clk, rst, out_s522, out_e522, result522);
PE P523(out_s491, out_e522, clk, rst, out_s523, out_e523, result523);
PE P524(out_s492, out_e523, clk, rst, out_s524, out_e524, result524);
PE P525(out_s493, out_e524, clk, rst, out_s525, out_e525, result525);
PE P526(out_s494, out_e525, clk, rst, out_s526, out_e526, result526);
PE P527(out_s495, out_e526, clk, rst, out_s527, out_e527, result527);
PE P528(out_s496, out_e527, clk, rst, out_s528, out_e528, result528);
PE P529(out_s497, out_e528, clk, rst, out_s529, out_e529, result529);
PE P530(out_s498, out_e529, clk, rst, out_s530, out_e530, result530);
PE P531(out_s499, out_e530, clk, rst, out_s531, out_e531, result531);
PE P532(out_s500, out_e531, clk, rst, out_s532, out_e532, result532);
PE P533(out_s501, out_e532, clk, rst, out_s533, out_e533, result533);
PE P534(out_s502, out_e533, clk, rst, out_s534, out_e534, result534);
PE P535(out_s503, out_e534, clk, rst, out_s535, out_e535, result535);
PE P536(out_s504, out_e535, clk, rst, out_s536, out_e536, result536);
PE P537(out_s505, out_e536, clk, rst, out_s537, out_e537, result537);
PE P538(out_s506, out_e537, clk, rst, out_s538, out_e538, result538);
PE P539(out_s507, out_e538, clk, rst, out_s539, out_e539, result539);
PE P540(out_s508, out_e539, clk, rst, out_s540, out_e540, result540);
PE P541(out_s509, out_e540, clk, rst, out_s541, out_e541, result541);
PE P542(out_s510, out_e541, clk, rst, out_s542, out_e542, result542);
PE P543(out_s511, out_e542, clk, rst, out_s543, out_e543, result543);

PE P545(out_s513, out_e544, clk, rst, out_s545, out_e545, result545);
PE P546(out_s514, out_e545, clk, rst, out_s546, out_e546, result546);
PE P547(out_s515, out_e546, clk, rst, out_s547, out_e547, result547);
PE P548(out_s516, out_e547, clk, rst, out_s548, out_e548, result548);
PE P549(out_s517, out_e548, clk, rst, out_s549, out_e549, result549);
PE P550(out_s518, out_e549, clk, rst, out_s550, out_e550, result550);
PE P551(out_s519, out_e550, clk, rst, out_s551, out_e551, result551);
PE P552(out_s520, out_e551, clk, rst, out_s552, out_e552, result552);
PE P553(out_s521, out_e552, clk, rst, out_s553, out_e553, result553);
PE P554(out_s522, out_e553, clk, rst, out_s554, out_e554, result554);
PE P555(out_s523, out_e554, clk, rst, out_s555, out_e555, result555);
PE P556(out_s524, out_e555, clk, rst, out_s556, out_e556, result556);
PE P557(out_s525, out_e556, clk, rst, out_s557, out_e557, result557);
PE P558(out_s526, out_e557, clk, rst, out_s558, out_e558, result558);
PE P559(out_s527, out_e558, clk, rst, out_s559, out_e559, result559);
PE P560(out_s528, out_e559, clk, rst, out_s560, out_e560, result560);
PE P561(out_s529, out_e560, clk, rst, out_s561, out_e561, result561);
PE P562(out_s530, out_e561, clk, rst, out_s562, out_e562, result562);
PE P563(out_s531, out_e562, clk, rst, out_s563, out_e563, result563);
PE P564(out_s532, out_e563, clk, rst, out_s564, out_e564, result564);
PE P565(out_s533, out_e564, clk, rst, out_s565, out_e565, result565);
PE P566(out_s534, out_e565, clk, rst, out_s566, out_e566, result566);
PE P567(out_s535, out_e566, clk, rst, out_s567, out_e567, result567);
PE P568(out_s536, out_e567, clk, rst, out_s568, out_e568, result568);
PE P569(out_s537, out_e568, clk, rst, out_s569, out_e569, result569);
PE P570(out_s538, out_e569, clk, rst, out_s570, out_e570, result570);
PE P571(out_s539, out_e570, clk, rst, out_s571, out_e571, result571);
PE P572(out_s540, out_e571, clk, rst, out_s572, out_e572, result572);
PE P573(out_s541, out_e572, clk, rst, out_s573, out_e573, result573);
PE P574(out_s542, out_e573, clk, rst, out_s574, out_e574, result574);
PE P575(out_s543, out_e574, clk, rst, out_s575, out_e575, result575);

PE P577(out_s545, out_e576, clk, rst, out_s577, out_e577, result577);
PE P578(out_s546, out_e577, clk, rst, out_s578, out_e578, result578);
PE P579(out_s547, out_e578, clk, rst, out_s579, out_e579, result579);
PE P580(out_s548, out_e579, clk, rst, out_s580, out_e580, result580);
PE P581(out_s549, out_e580, clk, rst, out_s581, out_e581, result581);
PE P582(out_s550, out_e581, clk, rst, out_s582, out_e582, result582);
PE P583(out_s551, out_e582, clk, rst, out_s583, out_e583, result583);
PE P584(out_s552, out_e583, clk, rst, out_s584, out_e584, result584);
PE P585(out_s553, out_e584, clk, rst, out_s585, out_e585, result585);
PE P586(out_s554, out_e585, clk, rst, out_s586, out_e586, result586);
PE P587(out_s555, out_e586, clk, rst, out_s587, out_e587, result587);
PE P588(out_s556, out_e587, clk, rst, out_s588, out_e588, result588);
PE P589(out_s557, out_e588, clk, rst, out_s589, out_e589, result589);
PE P590(out_s558, out_e589, clk, rst, out_s590, out_e590, result590);
PE P591(out_s559, out_e590, clk, rst, out_s591, out_e591, result591);
PE P592(out_s560, out_e591, clk, rst, out_s592, out_e592, result592);
PE P593(out_s561, out_e592, clk, rst, out_s593, out_e593, result593);
PE P594(out_s562, out_e593, clk, rst, out_s594, out_e594, result594);
PE P595(out_s563, out_e594, clk, rst, out_s595, out_e595, result595);
PE P596(out_s564, out_e595, clk, rst, out_s596, out_e596, result596);
PE P597(out_s565, out_e596, clk, rst, out_s597, out_e597, result597);
PE P598(out_s566, out_e597, clk, rst, out_s598, out_e598, result598);
PE P599(out_s567, out_e598, clk, rst, out_s599, out_e599, result599);
PE P600(out_s568, out_e599, clk, rst, out_s600, out_e600, result600);
PE P601(out_s569, out_e600, clk, rst, out_s601, out_e601, result601);
PE P602(out_s570, out_e601, clk, rst, out_s602, out_e602, result602);
PE P603(out_s571, out_e602, clk, rst, out_s603, out_e603, result603);
PE P604(out_s572, out_e603, clk, rst, out_s604, out_e604, result604);
PE P605(out_s573, out_e604, clk, rst, out_s605, out_e605, result605);
PE P606(out_s574, out_e605, clk, rst, out_s606, out_e606, result606);
PE P607(out_s575, out_e606, clk, rst, out_s607, out_e607, result607);

PE P609(out_s577, out_e608, clk, rst, out_s609, out_e609, result609);
PE P610(out_s578, out_e609, clk, rst, out_s610, out_e610, result610);
PE P611(out_s579, out_e610, clk, rst, out_s611, out_e611, result611);
PE P612(out_s580, out_e611, clk, rst, out_s612, out_e612, result612);
PE P613(out_s581, out_e612, clk, rst, out_s613, out_e613, result613);
PE P614(out_s582, out_e613, clk, rst, out_s614, out_e614, result614);
PE P615(out_s583, out_e614, clk, rst, out_s615, out_e615, result615);
PE P616(out_s584, out_e615, clk, rst, out_s616, out_e616, result616);
PE P617(out_s585, out_e616, clk, rst, out_s617, out_e617, result617);
PE P618(out_s586, out_e617, clk, rst, out_s618, out_e618, result618);
PE P619(out_s587, out_e618, clk, rst, out_s619, out_e619, result619);
PE P620(out_s588, out_e619, clk, rst, out_s620, out_e620, result620);
PE P621(out_s589, out_e620, clk, rst, out_s621, out_e621, result621);
PE P622(out_s590, out_e621, clk, rst, out_s622, out_e622, result622);
PE P623(out_s591, out_e622, clk, rst, out_s623, out_e623, result623);
PE P624(out_s592, out_e623, clk, rst, out_s624, out_e624, result624);
PE P625(out_s593, out_e624, clk, rst, out_s625, out_e625, result625);
PE P626(out_s594, out_e625, clk, rst, out_s626, out_e626, result626);
PE P627(out_s595, out_e626, clk, rst, out_s627, out_e627, result627);
PE P628(out_s596, out_e627, clk, rst, out_s628, out_e628, result628);
PE P629(out_s597, out_e628, clk, rst, out_s629, out_e629, result629);
PE P630(out_s598, out_e629, clk, rst, out_s630, out_e630, result630);
PE P631(out_s599, out_e630, clk, rst, out_s631, out_e631, result631);
PE P632(out_s600, out_e631, clk, rst, out_s632, out_e632, result632);
PE P633(out_s601, out_e632, clk, rst, out_s633, out_e633, result633);
PE P634(out_s602, out_e633, clk, rst, out_s634, out_e634, result634);
PE P635(out_s603, out_e634, clk, rst, out_s635, out_e635, result635);
PE P636(out_s604, out_e635, clk, rst, out_s636, out_e636, result636);
PE P637(out_s605, out_e636, clk, rst, out_s637, out_e637, result637);
PE P638(out_s606, out_e637, clk, rst, out_s638, out_e638, result638);
PE P639(out_s607, out_e638, clk, rst, out_s639, out_e639, result639);

PE P641(out_s609, out_e640, clk, rst, out_s641, out_e641, result641);
PE P642(out_s610, out_e641, clk, rst, out_s642, out_e642, result642);
PE P643(out_s611, out_e642, clk, rst, out_s643, out_e643, result643);
PE P644(out_s612, out_e643, clk, rst, out_s644, out_e644, result644);
PE P645(out_s613, out_e644, clk, rst, out_s645, out_e645, result645);
PE P646(out_s614, out_e645, clk, rst, out_s646, out_e646, result646);
PE P647(out_s615, out_e646, clk, rst, out_s647, out_e647, result647);
PE P648(out_s616, out_e647, clk, rst, out_s648, out_e648, result648);
PE P649(out_s617, out_e648, clk, rst, out_s649, out_e649, result649);
PE P650(out_s618, out_e649, clk, rst, out_s650, out_e650, result650);
PE P651(out_s619, out_e650, clk, rst, out_s651, out_e651, result651);
PE P652(out_s620, out_e651, clk, rst, out_s652, out_e652, result652);
PE P653(out_s621, out_e652, clk, rst, out_s653, out_e653, result653);
PE P654(out_s622, out_e653, clk, rst, out_s654, out_e654, result654);
PE P655(out_s623, out_e654, clk, rst, out_s655, out_e655, result655);
PE P656(out_s624, out_e655, clk, rst, out_s656, out_e656, result656);
PE P657(out_s625, out_e656, clk, rst, out_s657, out_e657, result657);
PE P658(out_s626, out_e657, clk, rst, out_s658, out_e658, result658);
PE P659(out_s627, out_e658, clk, rst, out_s659, out_e659, result659);
PE P660(out_s628, out_e659, clk, rst, out_s660, out_e660, result660);
PE P661(out_s629, out_e660, clk, rst, out_s661, out_e661, result661);
PE P662(out_s630, out_e661, clk, rst, out_s662, out_e662, result662);
PE P663(out_s631, out_e662, clk, rst, out_s663, out_e663, result663);
PE P664(out_s632, out_e663, clk, rst, out_s664, out_e664, result664);
PE P665(out_s633, out_e664, clk, rst, out_s665, out_e665, result665);
PE P666(out_s634, out_e665, clk, rst, out_s666, out_e666, result666);
PE P667(out_s635, out_e666, clk, rst, out_s667, out_e667, result667);
PE P668(out_s636, out_e667, clk, rst, out_s668, out_e668, result668);
PE P669(out_s637, out_e668, clk, rst, out_s669, out_e669, result669);
PE P670(out_s638, out_e669, clk, rst, out_s670, out_e670, result670);
PE P671(out_s639, out_e670, clk, rst, out_s671, out_e671, result671);

PE P673(out_s641, out_e672, clk, rst, out_s673, out_e673, result673);
PE P674(out_s642, out_e673, clk, rst, out_s674, out_e674, result674);
PE P675(out_s643, out_e674, clk, rst, out_s675, out_e675, result675);
PE P676(out_s644, out_e675, clk, rst, out_s676, out_e676, result676);
PE P677(out_s645, out_e676, clk, rst, out_s677, out_e677, result677);
PE P678(out_s646, out_e677, clk, rst, out_s678, out_e678, result678);
PE P679(out_s647, out_e678, clk, rst, out_s679, out_e679, result679);
PE P680(out_s648, out_e679, clk, rst, out_s680, out_e680, result680);
PE P681(out_s649, out_e680, clk, rst, out_s681, out_e681, result681);
PE P682(out_s650, out_e681, clk, rst, out_s682, out_e682, result682);
PE P683(out_s651, out_e682, clk, rst, out_s683, out_e683, result683);
PE P684(out_s652, out_e683, clk, rst, out_s684, out_e684, result684);
PE P685(out_s653, out_e684, clk, rst, out_s685, out_e685, result685);
PE P686(out_s654, out_e685, clk, rst, out_s686, out_e686, result686);
PE P687(out_s655, out_e686, clk, rst, out_s687, out_e687, result687);
PE P688(out_s656, out_e687, clk, rst, out_s688, out_e688, result688);
PE P689(out_s657, out_e688, clk, rst, out_s689, out_e689, result689);
PE P690(out_s658, out_e689, clk, rst, out_s690, out_e690, result690);
PE P691(out_s659, out_e690, clk, rst, out_s691, out_e691, result691);
PE P692(out_s660, out_e691, clk, rst, out_s692, out_e692, result692);
PE P693(out_s661, out_e692, clk, rst, out_s693, out_e693, result693);
PE P694(out_s662, out_e693, clk, rst, out_s694, out_e694, result694);
PE P695(out_s663, out_e694, clk, rst, out_s695, out_e695, result695);
PE P696(out_s664, out_e695, clk, rst, out_s696, out_e696, result696);
PE P697(out_s665, out_e696, clk, rst, out_s697, out_e697, result697);
PE P698(out_s666, out_e697, clk, rst, out_s698, out_e698, result698);
PE P699(out_s667, out_e698, clk, rst, out_s699, out_e699, result699);
PE P700(out_s668, out_e699, clk, rst, out_s700, out_e700, result700);
PE P701(out_s669, out_e700, clk, rst, out_s701, out_e701, result701);
PE P702(out_s670, out_e701, clk, rst, out_s702, out_e702, result702);
PE P703(out_s671, out_e702, clk, rst, out_s703, out_e703, result703);

PE P705(out_s673, out_e704, clk, rst, out_s705, out_e705, result705);
PE P706(out_s674, out_e705, clk, rst, out_s706, out_e706, result706);
PE P707(out_s675, out_e706, clk, rst, out_s707, out_e707, result707);
PE P708(out_s676, out_e707, clk, rst, out_s708, out_e708, result708);
PE P709(out_s677, out_e708, clk, rst, out_s709, out_e709, result709);
PE P710(out_s678, out_e709, clk, rst, out_s710, out_e710, result710);
PE P711(out_s679, out_e710, clk, rst, out_s711, out_e711, result711);
PE P712(out_s680, out_e711, clk, rst, out_s712, out_e712, result712);
PE P713(out_s681, out_e712, clk, rst, out_s713, out_e713, result713);
PE P714(out_s682, out_e713, clk, rst, out_s714, out_e714, result714);
PE P715(out_s683, out_e714, clk, rst, out_s715, out_e715, result715);
PE P716(out_s684, out_e715, clk, rst, out_s716, out_e716, result716);
PE P717(out_s685, out_e716, clk, rst, out_s717, out_e717, result717);
PE P718(out_s686, out_e717, clk, rst, out_s718, out_e718, result718);
PE P719(out_s687, out_e718, clk, rst, out_s719, out_e719, result719);
PE P720(out_s688, out_e719, clk, rst, out_s720, out_e720, result720);
PE P721(out_s689, out_e720, clk, rst, out_s721, out_e721, result721);
PE P722(out_s690, out_e721, clk, rst, out_s722, out_e722, result722);
PE P723(out_s691, out_e722, clk, rst, out_s723, out_e723, result723);
PE P724(out_s692, out_e723, clk, rst, out_s724, out_e724, result724);
PE P725(out_s693, out_e724, clk, rst, out_s725, out_e725, result725);
PE P726(out_s694, out_e725, clk, rst, out_s726, out_e726, result726);
PE P727(out_s695, out_e726, clk, rst, out_s727, out_e727, result727);
PE P728(out_s696, out_e727, clk, rst, out_s728, out_e728, result728);
PE P729(out_s697, out_e728, clk, rst, out_s729, out_e729, result729);
PE P730(out_s698, out_e729, clk, rst, out_s730, out_e730, result730);
PE P731(out_s699, out_e730, clk, rst, out_s731, out_e731, result731);
PE P732(out_s700, out_e731, clk, rst, out_s732, out_e732, result732);
PE P733(out_s701, out_e732, clk, rst, out_s733, out_e733, result733);
PE P734(out_s702, out_e733, clk, rst, out_s734, out_e734, result734);
PE P735(out_s703, out_e734, clk, rst, out_s735, out_e735, result735);

PE P737(out_s705, out_e736, clk, rst, out_s737, out_e737, result737);
PE P738(out_s706, out_e737, clk, rst, out_s738, out_e738, result738);
PE P739(out_s707, out_e738, clk, rst, out_s739, out_e739, result739);
PE P740(out_s708, out_e739, clk, rst, out_s740, out_e740, result740);
PE P741(out_s709, out_e740, clk, rst, out_s741, out_e741, result741);
PE P742(out_s710, out_e741, clk, rst, out_s742, out_e742, result742);
PE P743(out_s711, out_e742, clk, rst, out_s743, out_e743, result743);
PE P744(out_s712, out_e743, clk, rst, out_s744, out_e744, result744);
PE P745(out_s713, out_e744, clk, rst, out_s745, out_e745, result745);
PE P746(out_s714, out_e745, clk, rst, out_s746, out_e746, result746);
PE P747(out_s715, out_e746, clk, rst, out_s747, out_e747, result747);
PE P748(out_s716, out_e747, clk, rst, out_s748, out_e748, result748);
PE P749(out_s717, out_e748, clk, rst, out_s749, out_e749, result749);
PE P750(out_s718, out_e749, clk, rst, out_s750, out_e750, result750);
PE P751(out_s719, out_e750, clk, rst, out_s751, out_e751, result751);
PE P752(out_s720, out_e751, clk, rst, out_s752, out_e752, result752);
PE P753(out_s721, out_e752, clk, rst, out_s753, out_e753, result753);
PE P754(out_s722, out_e753, clk, rst, out_s754, out_e754, result754);
PE P755(out_s723, out_e754, clk, rst, out_s755, out_e755, result755);
PE P756(out_s724, out_e755, clk, rst, out_s756, out_e756, result756);
PE P757(out_s725, out_e756, clk, rst, out_s757, out_e757, result757);
PE P758(out_s726, out_e757, clk, rst, out_s758, out_e758, result758);
PE P759(out_s727, out_e758, clk, rst, out_s759, out_e759, result759);
PE P760(out_s728, out_e759, clk, rst, out_s760, out_e760, result760);
PE P761(out_s729, out_e760, clk, rst, out_s761, out_e761, result761);
PE P762(out_s730, out_e761, clk, rst, out_s762, out_e762, result762);
PE P763(out_s731, out_e762, clk, rst, out_s763, out_e763, result763);
PE P764(out_s732, out_e763, clk, rst, out_s764, out_e764, result764);
PE P765(out_s733, out_e764, clk, rst, out_s765, out_e765, result765);
PE P766(out_s734, out_e765, clk, rst, out_s766, out_e766, result766);
PE P767(out_s735, out_e766, clk, rst, out_s767, out_e767, result767);

PE P769(out_s737, out_e768, clk, rst, out_s769, out_e769, result769);
PE P770(out_s738, out_e769, clk, rst, out_s770, out_e770, result770);
PE P771(out_s739, out_e770, clk, rst, out_s771, out_e771, result771);
PE P772(out_s740, out_e771, clk, rst, out_s772, out_e772, result772);
PE P773(out_s741, out_e772, clk, rst, out_s773, out_e773, result773);
PE P774(out_s742, out_e773, clk, rst, out_s774, out_e774, result774);
PE P775(out_s743, out_e774, clk, rst, out_s775, out_e775, result775);
PE P776(out_s744, out_e775, clk, rst, out_s776, out_e776, result776);
PE P777(out_s745, out_e776, clk, rst, out_s777, out_e777, result777);
PE P778(out_s746, out_e777, clk, rst, out_s778, out_e778, result778);
PE P779(out_s747, out_e778, clk, rst, out_s779, out_e779, result779);
PE P780(out_s748, out_e779, clk, rst, out_s780, out_e780, result780);
PE P781(out_s749, out_e780, clk, rst, out_s781, out_e781, result781);
PE P782(out_s750, out_e781, clk, rst, out_s782, out_e782, result782);
PE P783(out_s751, out_e782, clk, rst, out_s783, out_e783, result783);
PE P784(out_s752, out_e783, clk, rst, out_s784, out_e784, result784);
PE P785(out_s753, out_e784, clk, rst, out_s785, out_e785, result785);
PE P786(out_s754, out_e785, clk, rst, out_s786, out_e786, result786);
PE P787(out_s755, out_e786, clk, rst, out_s787, out_e787, result787);
PE P788(out_s756, out_e787, clk, rst, out_s788, out_e788, result788);
PE P789(out_s757, out_e788, clk, rst, out_s789, out_e789, result789);
PE P790(out_s758, out_e789, clk, rst, out_s790, out_e790, result790);
PE P791(out_s759, out_e790, clk, rst, out_s791, out_e791, result791);
PE P792(out_s760, out_e791, clk, rst, out_s792, out_e792, result792);
PE P793(out_s761, out_e792, clk, rst, out_s793, out_e793, result793);
PE P794(out_s762, out_e793, clk, rst, out_s794, out_e794, result794);
PE P795(out_s763, out_e794, clk, rst, out_s795, out_e795, result795);
PE P796(out_s764, out_e795, clk, rst, out_s796, out_e796, result796);
PE P797(out_s765, out_e796, clk, rst, out_s797, out_e797, result797);
PE P798(out_s766, out_e797, clk, rst, out_s798, out_e798, result798);
PE P799(out_s767, out_e798, clk, rst, out_s799, out_e799, result799);

PE P801(out_s769, out_e800, clk, rst, out_s801, out_e801, result801);
PE P802(out_s770, out_e801, clk, rst, out_s802, out_e802, result802);
PE P803(out_s771, out_e802, clk, rst, out_s803, out_e803, result803);
PE P804(out_s772, out_e803, clk, rst, out_s804, out_e804, result804);
PE P805(out_s773, out_e804, clk, rst, out_s805, out_e805, result805);
PE P806(out_s774, out_e805, clk, rst, out_s806, out_e806, result806);
PE P807(out_s775, out_e806, clk, rst, out_s807, out_e807, result807);
PE P808(out_s776, out_e807, clk, rst, out_s808, out_e808, result808);
PE P809(out_s777, out_e808, clk, rst, out_s809, out_e809, result809);
PE P810(out_s778, out_e809, clk, rst, out_s810, out_e810, result810);
PE P811(out_s779, out_e810, clk, rst, out_s811, out_e811, result811);
PE P812(out_s780, out_e811, clk, rst, out_s812, out_e812, result812);
PE P813(out_s781, out_e812, clk, rst, out_s813, out_e813, result813);
PE P814(out_s782, out_e813, clk, rst, out_s814, out_e814, result814);
PE P815(out_s783, out_e814, clk, rst, out_s815, out_e815, result815);
PE P816(out_s784, out_e815, clk, rst, out_s816, out_e816, result816);
PE P817(out_s785, out_e816, clk, rst, out_s817, out_e817, result817);
PE P818(out_s786, out_e817, clk, rst, out_s818, out_e818, result818);
PE P819(out_s787, out_e818, clk, rst, out_s819, out_e819, result819);
PE P820(out_s788, out_e819, clk, rst, out_s820, out_e820, result820);
PE P821(out_s789, out_e820, clk, rst, out_s821, out_e821, result821);
PE P822(out_s790, out_e821, clk, rst, out_s822, out_e822, result822);
PE P823(out_s791, out_e822, clk, rst, out_s823, out_e823, result823);
PE P824(out_s792, out_e823, clk, rst, out_s824, out_e824, result824);
PE P825(out_s793, out_e824, clk, rst, out_s825, out_e825, result825);
PE P826(out_s794, out_e825, clk, rst, out_s826, out_e826, result826);
PE P827(out_s795, out_e826, clk, rst, out_s827, out_e827, result827);
PE P828(out_s796, out_e827, clk, rst, out_s828, out_e828, result828);
PE P829(out_s797, out_e828, clk, rst, out_s829, out_e829, result829);
PE P830(out_s798, out_e829, clk, rst, out_s830, out_e830, result830);
PE P831(out_s799, out_e830, clk, rst, out_s831, out_e831, result831);

PE P833(out_s801, out_e832, clk, rst, out_s833, out_e833, result833);
PE P834(out_s802, out_e833, clk, rst, out_s834, out_e834, result834);
PE P835(out_s803, out_e834, clk, rst, out_s835, out_e835, result835);
PE P836(out_s804, out_e835, clk, rst, out_s836, out_e836, result836);
PE P837(out_s805, out_e836, clk, rst, out_s837, out_e837, result837);
PE P838(out_s806, out_e837, clk, rst, out_s838, out_e838, result838);
PE P839(out_s807, out_e838, clk, rst, out_s839, out_e839, result839);
PE P840(out_s808, out_e839, clk, rst, out_s840, out_e840, result840);
PE P841(out_s809, out_e840, clk, rst, out_s841, out_e841, result841);
PE P842(out_s810, out_e841, clk, rst, out_s842, out_e842, result842);
PE P843(out_s811, out_e842, clk, rst, out_s843, out_e843, result843);
PE P844(out_s812, out_e843, clk, rst, out_s844, out_e844, result844);
PE P845(out_s813, out_e844, clk, rst, out_s845, out_e845, result845);
PE P846(out_s814, out_e845, clk, rst, out_s846, out_e846, result846);
PE P847(out_s815, out_e846, clk, rst, out_s847, out_e847, result847);
PE P848(out_s816, out_e847, clk, rst, out_s848, out_e848, result848);
PE P849(out_s817, out_e848, clk, rst, out_s849, out_e849, result849);
PE P850(out_s818, out_e849, clk, rst, out_s850, out_e850, result850);
PE P851(out_s819, out_e850, clk, rst, out_s851, out_e851, result851);
PE P852(out_s820, out_e851, clk, rst, out_s852, out_e852, result852);
PE P853(out_s821, out_e852, clk, rst, out_s853, out_e853, result853);
PE P854(out_s822, out_e853, clk, rst, out_s854, out_e854, result854);
PE P855(out_s823, out_e854, clk, rst, out_s855, out_e855, result855);
PE P856(out_s824, out_e855, clk, rst, out_s856, out_e856, result856);
PE P857(out_s825, out_e856, clk, rst, out_s857, out_e857, result857);
PE P858(out_s826, out_e857, clk, rst, out_s858, out_e858, result858);
PE P859(out_s827, out_e858, clk, rst, out_s859, out_e859, result859);
PE P860(out_s828, out_e859, clk, rst, out_s860, out_e860, result860);
PE P861(out_s829, out_e860, clk, rst, out_s861, out_e861, result861);
PE P862(out_s830, out_e861, clk, rst, out_s862, out_e862, result862);
PE P863(out_s831, out_e862, clk, rst, out_s863, out_e863, result863);

PE P865(out_s833, out_e864, clk, rst, out_s865, out_e865, result865);
PE P866(out_s834, out_e865, clk, rst, out_s866, out_e866, result866);
PE P867(out_s835, out_e866, clk, rst, out_s867, out_e867, result867);
PE P868(out_s836, out_e867, clk, rst, out_s868, out_e868, result868);
PE P869(out_s837, out_e868, clk, rst, out_s869, out_e869, result869);
PE P870(out_s838, out_e869, clk, rst, out_s870, out_e870, result870);
PE P871(out_s839, out_e870, clk, rst, out_s871, out_e871, result871);
PE P872(out_s840, out_e871, clk, rst, out_s872, out_e872, result872);
PE P873(out_s841, out_e872, clk, rst, out_s873, out_e873, result873);
PE P874(out_s842, out_e873, clk, rst, out_s874, out_e874, result874);
PE P875(out_s843, out_e874, clk, rst, out_s875, out_e875, result875);
PE P876(out_s844, out_e875, clk, rst, out_s876, out_e876, result876);
PE P877(out_s845, out_e876, clk, rst, out_s877, out_e877, result877);
PE P878(out_s846, out_e877, clk, rst, out_s878, out_e878, result878);
PE P879(out_s847, out_e878, clk, rst, out_s879, out_e879, result879);
PE P880(out_s848, out_e879, clk, rst, out_s880, out_e880, result880);
PE P881(out_s849, out_e880, clk, rst, out_s881, out_e881, result881);
PE P882(out_s850, out_e881, clk, rst, out_s882, out_e882, result882);
PE P883(out_s851, out_e882, clk, rst, out_s883, out_e883, result883);
PE P884(out_s852, out_e883, clk, rst, out_s884, out_e884, result884);
PE P885(out_s853, out_e884, clk, rst, out_s885, out_e885, result885);
PE P886(out_s854, out_e885, clk, rst, out_s886, out_e886, result886);
PE P887(out_s855, out_e886, clk, rst, out_s887, out_e887, result887);
PE P888(out_s856, out_e887, clk, rst, out_s888, out_e888, result888);
PE P889(out_s857, out_e888, clk, rst, out_s889, out_e889, result889);
PE P890(out_s858, out_e889, clk, rst, out_s890, out_e890, result890);
PE P891(out_s859, out_e890, clk, rst, out_s891, out_e891, result891);
PE P892(out_s860, out_e891, clk, rst, out_s892, out_e892, result892);
PE P893(out_s861, out_e892, clk, rst, out_s893, out_e893, result893);
PE P894(out_s862, out_e893, clk, rst, out_s894, out_e894, result894);
PE P895(out_s863, out_e894, clk, rst, out_s895, out_e895, result895);

PE P897(out_s865, out_e896, clk, rst, out_s897, out_e897, result897);
PE P898(out_s866, out_e897, clk, rst, out_s898, out_e898, result898);
PE P899(out_s867, out_e898, clk, rst, out_s899, out_e899, result899);
PE P900(out_s868, out_e899, clk, rst, out_s900, out_e900, result900);
PE P901(out_s869, out_e900, clk, rst, out_s901, out_e901, result901);
PE P902(out_s870, out_e901, clk, rst, out_s902, out_e902, result902);
PE P903(out_s871, out_e902, clk, rst, out_s903, out_e903, result903);
PE P904(out_s872, out_e903, clk, rst, out_s904, out_e904, result904);
PE P905(out_s873, out_e904, clk, rst, out_s905, out_e905, result905);
PE P906(out_s874, out_e905, clk, rst, out_s906, out_e906, result906);
PE P907(out_s875, out_e906, clk, rst, out_s907, out_e907, result907);
PE P908(out_s876, out_e907, clk, rst, out_s908, out_e908, result908);
PE P909(out_s877, out_e908, clk, rst, out_s909, out_e909, result909);
PE P910(out_s878, out_e909, clk, rst, out_s910, out_e910, result910);
PE P911(out_s879, out_e910, clk, rst, out_s911, out_e911, result911);
PE P912(out_s880, out_e911, clk, rst, out_s912, out_e912, result912);
PE P913(out_s881, out_e912, clk, rst, out_s913, out_e913, result913);
PE P914(out_s882, out_e913, clk, rst, out_s914, out_e914, result914);
PE P915(out_s883, out_e914, clk, rst, out_s915, out_e915, result915);
PE P916(out_s884, out_e915, clk, rst, out_s916, out_e916, result916);
PE P917(out_s885, out_e916, clk, rst, out_s917, out_e917, result917);
PE P918(out_s886, out_e917, clk, rst, out_s918, out_e918, result918);
PE P919(out_s887, out_e918, clk, rst, out_s919, out_e919, result919);
PE P920(out_s888, out_e919, clk, rst, out_s920, out_e920, result920);
PE P921(out_s889, out_e920, clk, rst, out_s921, out_e921, result921);
PE P922(out_s890, out_e921, clk, rst, out_s922, out_e922, result922);
PE P923(out_s891, out_e922, clk, rst, out_s923, out_e923, result923);
PE P924(out_s892, out_e923, clk, rst, out_s924, out_e924, result924);
PE P925(out_s893, out_e924, clk, rst, out_s925, out_e925, result925);
PE P926(out_s894, out_e925, clk, rst, out_s926, out_e926, result926);
PE P927(out_s895, out_e926, clk, rst, out_s927, out_e927, result927);

PE P929(out_s897, out_e928, clk, rst, out_s929, out_e929, result929);
PE P930(out_s898, out_e929, clk, rst, out_s930, out_e930, result930);
PE P931(out_s899, out_e930, clk, rst, out_s931, out_e931, result931);
PE P932(out_s900, out_e931, clk, rst, out_s932, out_e932, result932);
PE P933(out_s901, out_e932, clk, rst, out_s933, out_e933, result933);
PE P934(out_s902, out_e933, clk, rst, out_s934, out_e934, result934);
PE P935(out_s903, out_e934, clk, rst, out_s935, out_e935, result935);
PE P936(out_s904, out_e935, clk, rst, out_s936, out_e936, result936);
PE P937(out_s905, out_e936, clk, rst, out_s937, out_e937, result937);
PE P938(out_s906, out_e937, clk, rst, out_s938, out_e938, result938);
PE P939(out_s907, out_e938, clk, rst, out_s939, out_e939, result939);
PE P940(out_s908, out_e939, clk, rst, out_s940, out_e940, result940);
PE P941(out_s909, out_e940, clk, rst, out_s941, out_e941, result941);
PE P942(out_s910, out_e941, clk, rst, out_s942, out_e942, result942);
PE P943(out_s911, out_e942, clk, rst, out_s943, out_e943, result943);
PE P944(out_s912, out_e943, clk, rst, out_s944, out_e944, result944);
PE P945(out_s913, out_e944, clk, rst, out_s945, out_e945, result945);
PE P946(out_s914, out_e945, clk, rst, out_s946, out_e946, result946);
PE P947(out_s915, out_e946, clk, rst, out_s947, out_e947, result947);
PE P948(out_s916, out_e947, clk, rst, out_s948, out_e948, result948);
PE P949(out_s917, out_e948, clk, rst, out_s949, out_e949, result949);
PE P950(out_s918, out_e949, clk, rst, out_s950, out_e950, result950);
PE P951(out_s919, out_e950, clk, rst, out_s951, out_e951, result951);
PE P952(out_s920, out_e951, clk, rst, out_s952, out_e952, result952);
PE P953(out_s921, out_e952, clk, rst, out_s953, out_e953, result953);
PE P954(out_s922, out_e953, clk, rst, out_s954, out_e954, result954);
PE P955(out_s923, out_e954, clk, rst, out_s955, out_e955, result955);
PE P956(out_s924, out_e955, clk, rst, out_s956, out_e956, result956);
PE P957(out_s925, out_e956, clk, rst, out_s957, out_e957, result957);
PE P958(out_s926, out_e957, clk, rst, out_s958, out_e958, result958);
PE P959(out_s927, out_e958, clk, rst, out_s959, out_e959, result959);

PE P961(out_s929, out_e960, clk, rst, out_s961, out_e961, result961);
PE P962(out_s930, out_e961, clk, rst, out_s962, out_e962, result962);
PE P963(out_s931, out_e962, clk, rst, out_s963, out_e963, result963);
PE P964(out_s932, out_e963, clk, rst, out_s964, out_e964, result964);
PE P965(out_s933, out_e964, clk, rst, out_s965, out_e965, result965);
PE P966(out_s934, out_e965, clk, rst, out_s966, out_e966, result966);
PE P967(out_s935, out_e966, clk, rst, out_s967, out_e967, result967);
PE P968(out_s936, out_e967, clk, rst, out_s968, out_e968, result968);
PE P969(out_s937, out_e968, clk, rst, out_s969, out_e969, result969);
PE P970(out_s938, out_e969, clk, rst, out_s970, out_e970, result970);
PE P971(out_s939, out_e970, clk, rst, out_s971, out_e971, result971);
PE P972(out_s940, out_e971, clk, rst, out_s972, out_e972, result972);
PE P973(out_s941, out_e972, clk, rst, out_s973, out_e973, result973);
PE P974(out_s942, out_e973, clk, rst, out_s974, out_e974, result974);
PE P975(out_s943, out_e974, clk, rst, out_s975, out_e975, result975);
PE P976(out_s944, out_e975, clk, rst, out_s976, out_e976, result976);
PE P977(out_s945, out_e976, clk, rst, out_s977, out_e977, result977);
PE P978(out_s946, out_e977, clk, rst, out_s978, out_e978, result978);
PE P979(out_s947, out_e978, clk, rst, out_s979, out_e979, result979);
PE P980(out_s948, out_e979, clk, rst, out_s980, out_e980, result980);
PE P981(out_s949, out_e980, clk, rst, out_s981, out_e981, result981);
PE P982(out_s950, out_e981, clk, rst, out_s982, out_e982, result982);
PE P983(out_s951, out_e982, clk, rst, out_s983, out_e983, result983);
PE P984(out_s952, out_e983, clk, rst, out_s984, out_e984, result984);
PE P985(out_s953, out_e984, clk, rst, out_s985, out_e985, result985);
PE P986(out_s954, out_e985, clk, rst, out_s986, out_e986, result986);
PE P987(out_s955, out_e986, clk, rst, out_s987, out_e987, result987);
PE P988(out_s956, out_e987, clk, rst, out_s988, out_e988, result988);
PE P989(out_s957, out_e988, clk, rst, out_s989, out_e989, result989);
PE P990(out_s958, out_e989, clk, rst, out_s990, out_e990, result990);
PE P991(out_s959, out_e990, clk, rst, out_s991, out_e991, result991);

PE P993(out_s961, out_e992, clk, rst, out_s993, out_e993, result993);
PE P994(out_s962, out_e993, clk, rst, out_s994, out_e994, result994);
PE P995(out_s963, out_e994, clk, rst, out_s995, out_e995, result995);
PE P996(out_s964, out_e995, clk, rst, out_s996, out_e996, result996);
PE P997(out_s965, out_e996, clk, rst, out_s997, out_e997, result997);
PE P998(out_s966, out_e997, clk, rst, out_s998, out_e998, result998);
PE P999(out_s967, out_e998, clk, rst, out_s999, out_e999, result999);
PE P1000(out_s968, out_e999, clk, rst, out_s1000, out_e1000, result1000);
PE P1001(out_s969, out_e1000, clk, rst, out_s1001, out_e1001, result1001);
PE P1002(out_s970, out_e1001, clk, rst, out_s1002, out_e1002, result1002);
PE P1003(out_s971, out_e1002, clk, rst, out_s1003, out_e1003, result1003);
PE P1004(out_s972, out_e1003, clk, rst, out_s1004, out_e1004, result1004);
PE P1005(out_s973, out_e1004, clk, rst, out_s1005, out_e1005, result1005);
PE P1006(out_s974, out_e1005, clk, rst, out_s1006, out_e1006, result1006);
PE P1007(out_s975, out_e1006, clk, rst, out_s1007, out_e1007, result1007);
PE P1008(out_s976, out_e1007, clk, rst, out_s1008, out_e1008, result1008);
PE P1009(out_s977, out_e1008, clk, rst, out_s1009, out_e1009, result1009);
PE P1010(out_s978, out_e1009, clk, rst, out_s1010, out_e1010, result1010);
PE P1011(out_s979, out_e1010, clk, rst, out_s1011, out_e1011, result1011);
PE P1012(out_s980, out_e1011, clk, rst, out_s1012, out_e1012, result1012);
PE P1013(out_s981, out_e1012, clk, rst, out_s1013, out_e1013, result1013);
PE P1014(out_s982, out_e1013, clk, rst, out_s1014, out_e1014, result1014);
PE P1015(out_s983, out_e1014, clk, rst, out_s1015, out_e1015, result1015);
PE P1016(out_s984, out_e1015, clk, rst, out_s1016, out_e1016, result1016);
PE P1017(out_s985, out_e1016, clk, rst, out_s1017, out_e1017, result1017);
PE P1018(out_s986, out_e1017, clk, rst, out_s1018, out_e1018, result1018);
PE P1019(out_s987, out_e1018, clk, rst, out_s1019, out_e1019, result1019);
PE P1020(out_s988, out_e1019, clk, rst, out_s1020, out_e1020, result1020);
PE P1021(out_s989, out_e1020, clk, rst, out_s1021, out_e1021, result1021);
PE P1022(out_s990, out_e1021, clk, rst, out_s1022, out_e1022, result1022);
PE P1023(out_s991, out_e1022, clk, rst, out_s1023, out_e1023, result1023);

always @(posedge clk or posedge rst) begin
    if(rst) begin
        done <= 0;
        count <= 0;
    end
    else begin
		result_out0<=result0;
		result_out1<=result1;
		result_out2<=result2;
		result_out3<=result3;
		result_out4<=result4;
		result_out5<=result5;
		result_out6<=result6;
		result_out7<=result7;
		result_out8<=result8;
		result_out9<=result9;
		result_out10<=result10;
		result_out11<=result11;
		result_out12<=result12;
		result_out13<=result13;
		result_out14<=result14;
		result_out15<=result15;
		result_out16<=result16;
		result_out17<=result17;
		result_out18<=result18;
		result_out19<=result19;
		result_out20<=result20;
		result_out21<=result21;
		result_out22<=result22;
		result_out23<=result23;
		result_out24<=result24;
		result_out25<=result25;
		result_out26<=result26;
		result_out27<=result27;
		result_out28<=result28;
		result_out29<=result29;
		result_out30<=result30;
		result_out31<=result31;
		result_out32<=result32;
		result_out33<=result33;
		result_out34<=result34;
		result_out35<=result35;
		result_out36<=result36;
		result_out37<=result37;
		result_out38<=result38;
		result_out39<=result39;
		result_out40<=result40;
		result_out41<=result41;
		result_out42<=result42;
		result_out43<=result43;
		result_out44<=result44;
		result_out45<=result45;
		result_out46<=result46;
		result_out47<=result47;
		result_out48<=result48;
		result_out49<=result49;
		result_out50<=result50;
		result_out51<=result51;
		result_out52<=result52;
		result_out53<=result53;
		result_out54<=result54;
		result_out55<=result55;
		result_out56<=result56;
		result_out57<=result57;
		result_out58<=result58;
		result_out59<=result59;
		result_out60<=result60;
		result_out61<=result61;
		result_out62<=result62;
		result_out63<=result63;
		result_out64<=result64;
		result_out65<=result65;
		result_out66<=result66;
		result_out67<=result67;
		result_out68<=result68;
		result_out69<=result69;
		result_out70<=result70;
		result_out71<=result71;
		result_out72<=result72;
		result_out73<=result73;
		result_out74<=result74;
		result_out75<=result75;
		result_out76<=result76;
		result_out77<=result77;
		result_out78<=result78;
		result_out79<=result79;
		result_out80<=result80;
		result_out81<=result81;
		result_out82<=result82;
		result_out83<=result83;
		result_out84<=result84;
		result_out85<=result85;
		result_out86<=result86;
		result_out87<=result87;
		result_out88<=result88;
		result_out89<=result89;
		result_out90<=result90;
		result_out91<=result91;
		result_out92<=result92;
		result_out93<=result93;
		result_out94<=result94;
		result_out95<=result95;
		result_out96<=result96;
		result_out97<=result97;
		result_out98<=result98;
		result_out99<=result99;
		result_out100<=result100;
		result_out101<=result101;
		result_out102<=result102;
		result_out103<=result103;
		result_out104<=result104;
		result_out105<=result105;
		result_out106<=result106;
		result_out107<=result107;
		result_out108<=result108;
		result_out109<=result109;
		result_out110<=result110;
		result_out111<=result111;
		result_out112<=result112;
		result_out113<=result113;
		result_out114<=result114;
		result_out115<=result115;
		result_out116<=result116;
		result_out117<=result117;
		result_out118<=result118;
		result_out119<=result119;
		result_out120<=result120;
		result_out121<=result121;
		result_out122<=result122;
		result_out123<=result123;
		result_out124<=result124;
		result_out125<=result125;
		result_out126<=result126;
		result_out127<=result127;
		result_out128<=result128;
		result_out129<=result129;
		result_out130<=result130;
		result_out131<=result131;
		result_out132<=result132;
		result_out133<=result133;
		result_out134<=result134;
		result_out135<=result135;
		result_out136<=result136;
		result_out137<=result137;
		result_out138<=result138;
		result_out139<=result139;
		result_out140<=result140;
		result_out141<=result141;
		result_out142<=result142;
		result_out143<=result143;
		result_out144<=result144;
		result_out145<=result145;
		result_out146<=result146;
		result_out147<=result147;
		result_out148<=result148;
		result_out149<=result149;
		result_out150<=result150;
		result_out151<=result151;
		result_out152<=result152;
		result_out153<=result153;
		result_out154<=result154;
		result_out155<=result155;
		result_out156<=result156;
		result_out157<=result157;
		result_out158<=result158;
		result_out159<=result159;
		result_out160<=result160;
		result_out161<=result161;
		result_out162<=result162;
		result_out163<=result163;
		result_out164<=result164;
		result_out165<=result165;
		result_out166<=result166;
		result_out167<=result167;
		result_out168<=result168;
		result_out169<=result169;
		result_out170<=result170;
		result_out171<=result171;
		result_out172<=result172;
		result_out173<=result173;
		result_out174<=result174;
		result_out175<=result175;
		result_out176<=result176;
		result_out177<=result177;
		result_out178<=result178;
		result_out179<=result179;
		result_out180<=result180;
		result_out181<=result181;
		result_out182<=result182;
		result_out183<=result183;
		result_out184<=result184;
		result_out185<=result185;
		result_out186<=result186;
		result_out187<=result187;
		result_out188<=result188;
		result_out189<=result189;
		result_out190<=result190;
		result_out191<=result191;
		result_out192<=result192;
		result_out193<=result193;
		result_out194<=result194;
		result_out195<=result195;
		result_out196<=result196;
		result_out197<=result197;
		result_out198<=result198;
		result_out199<=result199;
		result_out200<=result200;
		result_out201<=result201;
		result_out202<=result202;
		result_out203<=result203;
		result_out204<=result204;
		result_out205<=result205;
		result_out206<=result206;
		result_out207<=result207;
		result_out208<=result208;
		result_out209<=result209;
		result_out210<=result210;
		result_out211<=result211;
		result_out212<=result212;
		result_out213<=result213;
		result_out214<=result214;
		result_out215<=result215;
		result_out216<=result216;
		result_out217<=result217;
		result_out218<=result218;
		result_out219<=result219;
		result_out220<=result220;
		result_out221<=result221;
		result_out222<=result222;
		result_out223<=result223;
		result_out224<=result224;
		result_out225<=result225;
		result_out226<=result226;
		result_out227<=result227;
		result_out228<=result228;
		result_out229<=result229;
		result_out230<=result230;
		result_out231<=result231;
		result_out232<=result232;
		result_out233<=result233;
		result_out234<=result234;
		result_out235<=result235;
		result_out236<=result236;
		result_out237<=result237;
		result_out238<=result238;
		result_out239<=result239;
		result_out240<=result240;
		result_out241<=result241;
		result_out242<=result242;
		result_out243<=result243;
		result_out244<=result244;
		result_out245<=result245;
		result_out246<=result246;
		result_out247<=result247;
		result_out248<=result248;
		result_out249<=result249;
		result_out250<=result250;
		result_out251<=result251;
		result_out252<=result252;
		result_out253<=result253;
		result_out254<=result254;
		result_out255<=result255;
		result_out256<=result256;
		result_out257<=result257;
		result_out258<=result258;
		result_out259<=result259;
		result_out260<=result260;
		result_out261<=result261;
		result_out262<=result262;
		result_out263<=result263;
		result_out264<=result264;
		result_out265<=result265;
		result_out266<=result266;
		result_out267<=result267;
		result_out268<=result268;
		result_out269<=result269;
		result_out270<=result270;
		result_out271<=result271;
		result_out272<=result272;
		result_out273<=result273;
		result_out274<=result274;
		result_out275<=result275;
		result_out276<=result276;
		result_out277<=result277;
		result_out278<=result278;
		result_out279<=result279;
		result_out280<=result280;
		result_out281<=result281;
		result_out282<=result282;
		result_out283<=result283;
		result_out284<=result284;
		result_out285<=result285;
		result_out286<=result286;
		result_out287<=result287;
		result_out288<=result288;
		result_out289<=result289;
		result_out290<=result290;
		result_out291<=result291;
		result_out292<=result292;
		result_out293<=result293;
		result_out294<=result294;
		result_out295<=result295;
		result_out296<=result296;
		result_out297<=result297;
		result_out298<=result298;
		result_out299<=result299;
		result_out300<=result300;
		result_out301<=result301;
		result_out302<=result302;
		result_out303<=result303;
		result_out304<=result304;
		result_out305<=result305;
		result_out306<=result306;
		result_out307<=result307;
		result_out308<=result308;
		result_out309<=result309;
		result_out310<=result310;
		result_out311<=result311;
		result_out312<=result312;
		result_out313<=result313;
		result_out314<=result314;
		result_out315<=result315;
		result_out316<=result316;
		result_out317<=result317;
		result_out318<=result318;
		result_out319<=result319;
		result_out320<=result320;
		result_out321<=result321;
		result_out322<=result322;
		result_out323<=result323;
		result_out324<=result324;
		result_out325<=result325;
		result_out326<=result326;
		result_out327<=result327;
		result_out328<=result328;
		result_out329<=result329;
		result_out330<=result330;
		result_out331<=result331;
		result_out332<=result332;
		result_out333<=result333;
		result_out334<=result334;
		result_out335<=result335;
		result_out336<=result336;
		result_out337<=result337;
		result_out338<=result338;
		result_out339<=result339;
		result_out340<=result340;
		result_out341<=result341;
		result_out342<=result342;
		result_out343<=result343;
		result_out344<=result344;
		result_out345<=result345;
		result_out346<=result346;
		result_out347<=result347;
		result_out348<=result348;
		result_out349<=result349;
		result_out350<=result350;
		result_out351<=result351;
		result_out352<=result352;
		result_out353<=result353;
		result_out354<=result354;
		result_out355<=result355;
		result_out356<=result356;
		result_out357<=result357;
		result_out358<=result358;
		result_out359<=result359;
		result_out360<=result360;
		result_out361<=result361;
		result_out362<=result362;
		result_out363<=result363;
		result_out364<=result364;
		result_out365<=result365;
		result_out366<=result366;
		result_out367<=result367;
		result_out368<=result368;
		result_out369<=result369;
		result_out370<=result370;
		result_out371<=result371;
		result_out372<=result372;
		result_out373<=result373;
		result_out374<=result374;
		result_out375<=result375;
		result_out376<=result376;
		result_out377<=result377;
		result_out378<=result378;
		result_out379<=result379;
		result_out380<=result380;
		result_out381<=result381;
		result_out382<=result382;
		result_out383<=result383;
		result_out384<=result384;
		result_out385<=result385;
		result_out386<=result386;
		result_out387<=result387;
		result_out388<=result388;
		result_out389<=result389;
		result_out390<=result390;
		result_out391<=result391;
		result_out392<=result392;
		result_out393<=result393;
		result_out394<=result394;
		result_out395<=result395;
		result_out396<=result396;
		result_out397<=result397;
		result_out398<=result398;
		result_out399<=result399;
		result_out400<=result400;
		result_out401<=result401;
		result_out402<=result402;
		result_out403<=result403;
		result_out404<=result404;
		result_out405<=result405;
		result_out406<=result406;
		result_out407<=result407;
		result_out408<=result408;
		result_out409<=result409;
		result_out410<=result410;
		result_out411<=result411;
		result_out412<=result412;
		result_out413<=result413;
		result_out414<=result414;
		result_out415<=result415;
		result_out416<=result416;
		result_out417<=result417;
		result_out418<=result418;
		result_out419<=result419;
		result_out420<=result420;
		result_out421<=result421;
		result_out422<=result422;
		result_out423<=result423;
		result_out424<=result424;
		result_out425<=result425;
		result_out426<=result426;
		result_out427<=result427;
		result_out428<=result428;
		result_out429<=result429;
		result_out430<=result430;
		result_out431<=result431;
		result_out432<=result432;
		result_out433<=result433;
		result_out434<=result434;
		result_out435<=result435;
		result_out436<=result436;
		result_out437<=result437;
		result_out438<=result438;
		result_out439<=result439;
		result_out440<=result440;
		result_out441<=result441;
		result_out442<=result442;
		result_out443<=result443;
		result_out444<=result444;
		result_out445<=result445;
		result_out446<=result446;
		result_out447<=result447;
		result_out448<=result448;
		result_out449<=result449;
		result_out450<=result450;
		result_out451<=result451;
		result_out452<=result452;
		result_out453<=result453;
		result_out454<=result454;
		result_out455<=result455;
		result_out456<=result456;
		result_out457<=result457;
		result_out458<=result458;
		result_out459<=result459;
		result_out460<=result460;
		result_out461<=result461;
		result_out462<=result462;
		result_out463<=result463;
		result_out464<=result464;
		result_out465<=result465;
		result_out466<=result466;
		result_out467<=result467;
		result_out468<=result468;
		result_out469<=result469;
		result_out470<=result470;
		result_out471<=result471;
		result_out472<=result472;
		result_out473<=result473;
		result_out474<=result474;
		result_out475<=result475;
		result_out476<=result476;
		result_out477<=result477;
		result_out478<=result478;
		result_out479<=result479;
		result_out480<=result480;
		result_out481<=result481;
		result_out482<=result482;
		result_out483<=result483;
		result_out484<=result484;
		result_out485<=result485;
		result_out486<=result486;
		result_out487<=result487;
		result_out488<=result488;
		result_out489<=result489;
		result_out490<=result490;
		result_out491<=result491;
		result_out492<=result492;
		result_out493<=result493;
		result_out494<=result494;
		result_out495<=result495;
		result_out496<=result496;
		result_out497<=result497;
		result_out498<=result498;
		result_out499<=result499;
		result_out500<=result500;
		result_out501<=result501;
		result_out502<=result502;
		result_out503<=result503;
		result_out504<=result504;
		result_out505<=result505;
		result_out506<=result506;
		result_out507<=result507;
		result_out508<=result508;
		result_out509<=result509;
		result_out510<=result510;
		result_out511<=result511;
		result_out512<=result512;
		result_out513<=result513;
		result_out514<=result514;
		result_out515<=result515;
		result_out516<=result516;
		result_out517<=result517;
		result_out518<=result518;
		result_out519<=result519;
		result_out520<=result520;
		result_out521<=result521;
		result_out522<=result522;
		result_out523<=result523;
		result_out524<=result524;
		result_out525<=result525;
		result_out526<=result526;
		result_out527<=result527;
		result_out528<=result528;
		result_out529<=result529;
		result_out530<=result530;
		result_out531<=result531;
		result_out532<=result532;
		result_out533<=result533;
		result_out534<=result534;
		result_out535<=result535;
		result_out536<=result536;
		result_out537<=result537;
		result_out538<=result538;
		result_out539<=result539;
		result_out540<=result540;
		result_out541<=result541;
		result_out542<=result542;
		result_out543<=result543;
		result_out544<=result544;
		result_out545<=result545;
		result_out546<=result546;
		result_out547<=result547;
		result_out548<=result548;
		result_out549<=result549;
		result_out550<=result550;
		result_out551<=result551;
		result_out552<=result552;
		result_out553<=result553;
		result_out554<=result554;
		result_out555<=result555;
		result_out556<=result556;
		result_out557<=result557;
		result_out558<=result558;
		result_out559<=result559;
		result_out560<=result560;
		result_out561<=result561;
		result_out562<=result562;
		result_out563<=result563;
		result_out564<=result564;
		result_out565<=result565;
		result_out566<=result566;
		result_out567<=result567;
		result_out568<=result568;
		result_out569<=result569;
		result_out570<=result570;
		result_out571<=result571;
		result_out572<=result572;
		result_out573<=result573;
		result_out574<=result574;
		result_out575<=result575;
		result_out576<=result576;
		result_out577<=result577;
		result_out578<=result578;
		result_out579<=result579;
		result_out580<=result580;
		result_out581<=result581;
		result_out582<=result582;
		result_out583<=result583;
		result_out584<=result584;
		result_out585<=result585;
		result_out586<=result586;
		result_out587<=result587;
		result_out588<=result588;
		result_out589<=result589;
		result_out590<=result590;
		result_out591<=result591;
		result_out592<=result592;
		result_out593<=result593;
		result_out594<=result594;
		result_out595<=result595;
		result_out596<=result596;
		result_out597<=result597;
		result_out598<=result598;
		result_out599<=result599;
		result_out600<=result600;
		result_out601<=result601;
		result_out602<=result602;
		result_out603<=result603;
		result_out604<=result604;
		result_out605<=result605;
		result_out606<=result606;
		result_out607<=result607;
		result_out608<=result608;
		result_out609<=result609;
		result_out610<=result610;
		result_out611<=result611;
		result_out612<=result612;
		result_out613<=result613;
		result_out614<=result614;
		result_out615<=result615;
		result_out616<=result616;
		result_out617<=result617;
		result_out618<=result618;
		result_out619<=result619;
		result_out620<=result620;
		result_out621<=result621;
		result_out622<=result622;
		result_out623<=result623;
		result_out624<=result624;
		result_out625<=result625;
		result_out626<=result626;
		result_out627<=result627;
		result_out628<=result628;
		result_out629<=result629;
		result_out630<=result630;
		result_out631<=result631;
		result_out632<=result632;
		result_out633<=result633;
		result_out634<=result634;
		result_out635<=result635;
		result_out636<=result636;
		result_out637<=result637;
		result_out638<=result638;
		result_out639<=result639;
		result_out640<=result640;
		result_out641<=result641;
		result_out642<=result642;
		result_out643<=result643;
		result_out644<=result644;
		result_out645<=result645;
		result_out646<=result646;
		result_out647<=result647;
		result_out648<=result648;
		result_out649<=result649;
		result_out650<=result650;
		result_out651<=result651;
		result_out652<=result652;
		result_out653<=result653;
		result_out654<=result654;
		result_out655<=result655;
		result_out656<=result656;
		result_out657<=result657;
		result_out658<=result658;
		result_out659<=result659;
		result_out660<=result660;
		result_out661<=result661;
		result_out662<=result662;
		result_out663<=result663;
		result_out664<=result664;
		result_out665<=result665;
		result_out666<=result666;
		result_out667<=result667;
		result_out668<=result668;
		result_out669<=result669;
		result_out670<=result670;
		result_out671<=result671;
		result_out672<=result672;
		result_out673<=result673;
		result_out674<=result674;
		result_out675<=result675;
		result_out676<=result676;
		result_out677<=result677;
		result_out678<=result678;
		result_out679<=result679;
		result_out680<=result680;
		result_out681<=result681;
		result_out682<=result682;
		result_out683<=result683;
		result_out684<=result684;
		result_out685<=result685;
		result_out686<=result686;
		result_out687<=result687;
		result_out688<=result688;
		result_out689<=result689;
		result_out690<=result690;
		result_out691<=result691;
		result_out692<=result692;
		result_out693<=result693;
		result_out694<=result694;
		result_out695<=result695;
		result_out696<=result696;
		result_out697<=result697;
		result_out698<=result698;
		result_out699<=result699;
		result_out700<=result700;
		result_out701<=result701;
		result_out702<=result702;
		result_out703<=result703;
		result_out704<=result704;
		result_out705<=result705;
		result_out706<=result706;
		result_out707<=result707;
		result_out708<=result708;
		result_out709<=result709;
		result_out710<=result710;
		result_out711<=result711;
		result_out712<=result712;
		result_out713<=result713;
		result_out714<=result714;
		result_out715<=result715;
		result_out716<=result716;
		result_out717<=result717;
		result_out718<=result718;
		result_out719<=result719;
		result_out720<=result720;
		result_out721<=result721;
		result_out722<=result722;
		result_out723<=result723;
		result_out724<=result724;
		result_out725<=result725;
		result_out726<=result726;
		result_out727<=result727;
		result_out728<=result728;
		result_out729<=result729;
		result_out730<=result730;
		result_out731<=result731;
		result_out732<=result732;
		result_out733<=result733;
		result_out734<=result734;
		result_out735<=result735;
		result_out736<=result736;
		result_out737<=result737;
		result_out738<=result738;
		result_out739<=result739;
		result_out740<=result740;
		result_out741<=result741;
		result_out742<=result742;
		result_out743<=result743;
		result_out744<=result744;
		result_out745<=result745;
		result_out746<=result746;
		result_out747<=result747;
		result_out748<=result748;
		result_out749<=result749;
		result_out750<=result750;
		result_out751<=result751;
		result_out752<=result752;
		result_out753<=result753;
		result_out754<=result754;
		result_out755<=result755;
		result_out756<=result756;
		result_out757<=result757;
		result_out758<=result758;
		result_out759<=result759;
		result_out760<=result760;
		result_out761<=result761;
		result_out762<=result762;
		result_out763<=result763;
		result_out764<=result764;
		result_out765<=result765;
		result_out766<=result766;
		result_out767<=result767;
		result_out768<=result768;
		result_out769<=result769;
		result_out770<=result770;
		result_out771<=result771;
		result_out772<=result772;
		result_out773<=result773;
		result_out774<=result774;
		result_out775<=result775;
		result_out776<=result776;
		result_out777<=result777;
		result_out778<=result778;
		result_out779<=result779;
		result_out780<=result780;
		result_out781<=result781;
		result_out782<=result782;
		result_out783<=result783;
		result_out784<=result784;
		result_out785<=result785;
		result_out786<=result786;
		result_out787<=result787;
		result_out788<=result788;
		result_out789<=result789;
		result_out790<=result790;
		result_out791<=result791;
		result_out792<=result792;
		result_out793<=result793;
		result_out794<=result794;
		result_out795<=result795;
		result_out796<=result796;
		result_out797<=result797;
		result_out798<=result798;
		result_out799<=result799;
		result_out800<=result800;
		result_out801<=result801;
		result_out802<=result802;
		result_out803<=result803;
		result_out804<=result804;
		result_out805<=result805;
		result_out806<=result806;
		result_out807<=result807;
		result_out808<=result808;
		result_out809<=result809;
		result_out810<=result810;
		result_out811<=result811;
		result_out812<=result812;
		result_out813<=result813;
		result_out814<=result814;
		result_out815<=result815;
		result_out816<=result816;
		result_out817<=result817;
		result_out818<=result818;
		result_out819<=result819;
		result_out820<=result820;
		result_out821<=result821;
		result_out822<=result822;
		result_out823<=result823;
		result_out824<=result824;
		result_out825<=result825;
		result_out826<=result826;
		result_out827<=result827;
		result_out828<=result828;
		result_out829<=result829;
		result_out830<=result830;
		result_out831<=result831;
		result_out832<=result832;
		result_out833<=result833;
		result_out834<=result834;
		result_out835<=result835;
		result_out836<=result836;
		result_out837<=result837;
		result_out838<=result838;
		result_out839<=result839;
		result_out840<=result840;
		result_out841<=result841;
		result_out842<=result842;
		result_out843<=result843;
		result_out844<=result844;
		result_out845<=result845;
		result_out846<=result846;
		result_out847<=result847;
		result_out848<=result848;
		result_out849<=result849;
		result_out850<=result850;
		result_out851<=result851;
		result_out852<=result852;
		result_out853<=result853;
		result_out854<=result854;
		result_out855<=result855;
		result_out856<=result856;
		result_out857<=result857;
		result_out858<=result858;
		result_out859<=result859;
		result_out860<=result860;
		result_out861<=result861;
		result_out862<=result862;
		result_out863<=result863;
		result_out864<=result864;
		result_out865<=result865;
		result_out866<=result866;
		result_out867<=result867;
		result_out868<=result868;
		result_out869<=result869;
		result_out870<=result870;
		result_out871<=result871;
		result_out872<=result872;
		result_out873<=result873;
		result_out874<=result874;
		result_out875<=result875;
		result_out876<=result876;
		result_out877<=result877;
		result_out878<=result878;
		result_out879<=result879;
		result_out880<=result880;
		result_out881<=result881;
		result_out882<=result882;
		result_out883<=result883;
		result_out884<=result884;
		result_out885<=result885;
		result_out886<=result886;
		result_out887<=result887;
		result_out888<=result888;
		result_out889<=result889;
		result_out890<=result890;
		result_out891<=result891;
		result_out892<=result892;
		result_out893<=result893;
		result_out894<=result894;
		result_out895<=result895;
		result_out896<=result896;
		result_out897<=result897;
		result_out898<=result898;
		result_out899<=result899;
		result_out900<=result900;
		result_out901<=result901;
		result_out902<=result902;
		result_out903<=result903;
		result_out904<=result904;
		result_out905<=result905;
		result_out906<=result906;
		result_out907<=result907;
		result_out908<=result908;
		result_out909<=result909;
		result_out910<=result910;
		result_out911<=result911;
		result_out912<=result912;
		result_out913<=result913;
		result_out914<=result914;
		result_out915<=result915;
		result_out916<=result916;
		result_out917<=result917;
		result_out918<=result918;
		result_out919<=result919;
		result_out920<=result920;
		result_out921<=result921;
		result_out922<=result922;
		result_out923<=result923;
		result_out924<=result924;
		result_out925<=result925;
		result_out926<=result926;
		result_out927<=result927;
		result_out928<=result928;
		result_out929<=result929;
		result_out930<=result930;
		result_out931<=result931;
		result_out932<=result932;
		result_out933<=result933;
		result_out934<=result934;
		result_out935<=result935;
		result_out936<=result936;
		result_out937<=result937;
		result_out938<=result938;
		result_out939<=result939;
		result_out940<=result940;
		result_out941<=result941;
		result_out942<=result942;
		result_out943<=result943;
		result_out944<=result944;
		result_out945<=result945;
		result_out946<=result946;
		result_out947<=result947;
		result_out948<=result948;
		result_out949<=result949;
		result_out950<=result950;
		result_out951<=result951;
		result_out952<=result952;
		result_out953<=result953;
		result_out954<=result954;
		result_out955<=result955;
		result_out956<=result956;
		result_out957<=result957;
		result_out958<=result958;
		result_out959<=result959;
		result_out960<=result960;
		result_out961<=result961;
		result_out962<=result962;
		result_out963<=result963;
		result_out964<=result964;
		result_out965<=result965;
		result_out966<=result966;
		result_out967<=result967;
		result_out968<=result968;
		result_out969<=result969;
		result_out970<=result970;
		result_out971<=result971;
		result_out972<=result972;
		result_out973<=result973;
		result_out974<=result974;
		result_out975<=result975;
		result_out976<=result976;
		result_out977<=result977;
		result_out978<=result978;
		result_out979<=result979;
		result_out980<=result980;
		result_out981<=result981;
		result_out982<=result982;
		result_out983<=result983;
		result_out984<=result984;
		result_out985<=result985;
		result_out986<=result986;
		result_out987<=result987;
		result_out988<=result988;
		result_out989<=result989;
		result_out990<=result990;
		result_out991<=result991;
		result_out992<=result992;
		result_out993<=result993;
		result_out994<=result994;
		result_out995<=result995;
		result_out996<=result996;
		result_out997<=result997;
		result_out998<=result998;
		result_out999<=result999;
		result_out1000<=result1000;
		result_out1001<=result1001;
		result_out1002<=result1002;
		result_out1003<=result1003;
		result_out1004<=result1004;
		result_out1005<=result1005;
		result_out1006<=result1006;
		result_out1007<=result1007;
		result_out1008<=result1008;
		result_out1009<=result1009;
		result_out1010<=result1010;
		result_out1011<=result1011;
		result_out1012<=result1012;
		result_out1013<=result1013;
		result_out1014<=result1014;
		result_out1015<=result1015;
		result_out1016<=result1016;
		result_out1017<=result1017;
		result_out1018<=result1018;
		result_out1019<=result1019;
		result_out1020<=result1020;
		result_out1021<=result1021;
		result_out1022<=result1022;
		result_out1023<=result1023;
		if(count == 94) begin
            done <= 1;
            count <= 0;
        end
        else begin
            done <= 0;
            count <= count + 1;
        end
    end
end
endmodule
